��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F�)	�ŀ)v�ޑ"^��F��L�> Ó�����M4G�h�.Yv~��f�+�E�9�?���;�Ω0�4��H�;uS%."q��Zd�/�]�+G|��Ԇբ�n�<!�?�a,��5_��=�n�����~t��^}��ٸ�/��eLУvi�i���m�ޮ%G����i�}	�71\&��cq����+�zE��<�`\�L^�e�|�ی�k��=OV�B�v�@�1�^'盾�R��9��'E�򛚤�p�E^΂�Ok��������aG|#�	[m���}�����R��=��ئ4�r-����[�}�x� �|�LW!�c\j��:���ȳ�oi����_v����jqQ�#�d^��Fџ��<0�
)ߪw�B��ֺo\�s)��M�[��	�h_*9o��E_���]��F~�#?ٌp�&�5d1�)G+��� �n���?z!H��x8��U2�#��#T�I�%j=�մ� �Q��9n��C�)��Y���h2�'����lw��9\7�� �9�`�ꌗe��c^E���2;�%�R��� �w�Pk����9���sr~P����u|&��S�-�}	%N��v��	T)%O̘z#i!_ ���*�w�3�Ļ4�L�~�Ǌ���R�o��%!��V��R�����	+ښu�u��a� b� �$ɓ���������G��*�N�
?A}��02��߫w�<s�O������!&v��šc�lA��&���h�"@$��H��r�l�f)��b8�ۘ7c ���|�(<�1��Yh������*�㋽.L��E0pa'E���d�0E�J���G�?�X��$�fxo�#5�P}����,����w��g�VN�V
�#HȎ��U���̏��;Y��c4�p�C��Y9�\v	�5�MX��Ǌ��%�1��9x��X���Zk���j2 �5)e�-oO�P�]�ѐ��n���F�T����
)�@�s��t�P�܆�,\F�Ehi1�������"W�_e�y�ͦ�>>~�/��};�Ӈ�1�GҢ�m�����
 \ n���&��z��e��� ԺU��欀�Iv�˴��D�}!Kdh@����q(6ڮ��X�J&n��$�wݣY�=^'�1/NΖ�o�y�:ϱ���Ï
IL��i$����AI�
�g��i({w)�9��"畠��������dA`��=R�i)��}2"Tm$l)�2ٽ}ɷCf�&�y�K�E���Hi>���z,��ހZ�SqQ��ۘhyZ/��8��'v_JR�~jw1���n����g���{qE��8a��SE�o�u榩������6Y���R���m�{tA�!��N*N�zk��������n�UYy�W����L�����#�w��3�A�R��̮�KsU�H����U_�وo�d�n�1��t&%��U��D G�W/$Rh	�Ƨ��oQhM�6�w��1,�B!|�o���XO[�&�G[:�F�1:���3����ΐʴ��_76Q֋{s����۱�c_�O9j!�4��:����:l��U1y�J�Cм�6����5j�bf�	�fu�i��}yP�2֜:�~��	��Aw@�TeJ�*	��UyG5��Xz����	aby	J�)*��L{?0��s�BO��D�c�2�)�A��W7a�E��} �<�=�p�W�X- t,�k�yT4<dN�R�
x��3Ŭ����h�1!��j��]&��U"��f*�ڎxA���~�J9��~�kfn�W"�!J#D�����u����M�F�.�Q�M� /���)Dn1�;�Hw�'�?Y'��w�������'���\�BW��B��60��;�3<�{9���s��sg�b���pgpPk��a�Y[���#ʔ9��(��W핃��izh+��+���V�W"�`�-{�%��F�sTR�)����f�e�Z�.?���¡GVG��YH�ܣ����p� ��=k�;y���í�x���ȇ�?��Y1na��2s�cZ3^���{1���O��]`?�W	ʽ�x#VʍQ������z�M��&.sib�Z0O	�3��~��߽-���}��=�=�S����`U��O1�$��9��1�������|*v;��aD�ڳ�����Шvdb�ț���i>�xଆ�X|[0�,LI�)ˌZ�����]��e���t�_�kvf;iP��摴��Ǘ�
�@@��F����?e"ݬֻ��n�Q�F�'G��O���� W��a*������f�"��8Ŷ�p�W.�`�0��ya`�r�|ֲ��2<R�:%�i�cb�:5���4F�Sv[�ʫeq�~5�|�I) ���l|9���뛀G����Ϳ�x�\1�
��N�j��^
H|���=�}�H��X�(�=��N<!��,7��Vu��������	F�#k9�p2�4R~��:�%e0�@6�y��.�[����|%q�Hթ:����]�w�, ��l_�N��P.s�n�/�S�B��<���h�=�iu�p�RL��4�n���6��.)���1�-�^]�*v����p�R�;~�Ad��K1=rM�����4c/�tc�Ò2\ęD�C�k�.���֦�9@��o��VǑ�|�_]$(������$FA@XKS�m+���t�Y'�ߥF�甁~�)[�~�Bm,��� �콼/	��{��&��xɶ\
�4
jZ�F��`�E���*}����e$ T6+���#hMu��h|5|�1�L�U�>h,�"�޲�{��g�w.^�X\/�� P
O.�Yg��C� +C}p�
�kp���|K�6��A��q6���^��޾hAn�OC�G���>���2إ�J�J+�ǿ?-��h94��L�%����c�ͺ(R���]�]�Q���0sc�sտe���I�$F�TeL��>�/��ӣ�IpX���g����R�t����eA:m�a�n)�Q}l'(�^s���VҔ-3EC�Bu�"��5���]BW`t�iQb�	��0w���J9ǛK6e-L���n�7�w���C/c8��@��ު%:�t���a�1���WQr��A�kb����\K�0�Y }�q��?��������>W�C[�-���nh� v��$�kt��v��Ym����lRh�?�/%�im�_�8?E!��%w�]A۱�9�~|;�� �����iZ�,C�X������М�W'�.;�7�������z[�|��r�B}�ǈA�V/ǰ�M:	2���� ��I��piKlI��S4f�� �"���=�>����hj�t��K���xx��L��ko@^�U�ܛ���~���9GF�t�j*ŵ84���Uodp"D��X�Cxɞ>Ql��8�zI��ƿ���x'��^H2���2�X���)�����i��#�7��>H��~���)
P0��h�؄�z"Y�s�ݕGxw���g�yc�X��ͣ$�,'ڍp�V��zRg_J(�!�3{~5��O��D�
�٠��-���P�Dl�����}t�y8Mw޼)��N(l�\�����,~�<EHW��-�(!�a_)FA���i�
2�����P:/i�n��Dd�%�7��\6������W�#F՘քD�y���}�Ka�O�����Mz���O����h �Vn�W���9
������ x(����<����|?������`Z�&8�X�<�V�l����Ν֗�؜��r�g��@e⩉zUI����Tw*>;���3b��;+|;b�UNE� ��APN��)���Xa�9�5Dֽ
vEV������ ������Qm�qι���qU�h���@�����<��cQK���Vj+-[��� � <6Q�K�ω'=P�p�G
PB�E�r�x��o���4��K�ű���? W"�/H4|�w6�KC�ǰj7��ڜȵ(���w��%�����c��8
���w��F��������p�T�(���*=s��ٌ����ӇH8{�"o%'�Uf��@�̣����.CE`�V�@���K��Jo�@0+��%2�}#dف�{��]	8JDnj,����l��{�2,86�z58x
&N4������|��$þA���+�����Xe���6$�P��8T��6�X�{R��h3űi�bj_�T6�gÑ�H���p�r���^�㫼��L��@W2�W�T��
"8�H����~h��x#�aNf���!�����]���@zg��@�puF�5XN-	��!R߁wKb8�T+���MX�$� ��SJkG��w!H�=[?�� �cqc��^��:����?.50ߥF&���Q�I�u�X�Yj�g���G)���Y��hҝ%q����ܯ�t����%�O:|��И}"��Pb=N�,�n@1Ex��8C1�F6��|�(;\��kL�9C��B�)�+���mkҞX/�t��5�ҝTf�jA�2����D����i�o�:B��ƶ���~t:�O�@�9j_A�_���591 �51o��nip{3����M����]ɹR�	���6WR/5��F5�W�8*����"�,��6V��Z	�R�2>�"�\U�K�(��E��o��4jP��X"�i�):d�hqU�>���O��r�F�\��Sf��Y�`�S
Z��C�n��DB.�����?���|V�_�� p���!�7��B���O�x��}W����-��:�p�K6�������0�	�6�.���\���$��Bb���sߩ�-	W��*��:l�zн��Zy�x/�A�W���O�RgW�91��%7M�̮�M�BE�'�8��Y0&�@5﨓��b�T��+!Rw�}�æ9��Z2v��ٺ)�p����R;_I���鼉�������0j������3�2%/�Q$���	Q�)�IƬQ��InZ� �Ј�A&G��q�ɹo��&v�0v�Dmw��X�E��&�i�vT_?�VNW%E�]��Tʊ��I���!���;�:����c�G�D��Јx�n��re&����cLm*���P9��1��RV)��hڶ�����"��xHW)ެ��G]b�S�$Y0��5)���=�av�~��S�:r}+_�C&��*_��!w-O�"u��&g�JW'L�2`5���	��ӽZQv�©%������ 4.�Xznd?H��踉n�o�}udz��E#_�	]"��ju���R�卹�ހ$�V�iv�gyN�珱@��g���h�`�#I�������-���������co���&O�I���3�Y
�!�y)r�X����c�W�ᢁ���x{p��[?o�˗�9OA:�X�8%O)XZ���K�p�L�bH��j�۷!ŕ�&�B|�F�f#�mśE�r��`��dR�s��9�kK�F;2;�7�8׬�v~�#F �=�1�$��UӇ�(�I������a]Q���T������!w:�9g�n�z�-�w}}�<�$��_^��_ЮM4qA��f�Ϧ�$q�u�Ġ��Оˬ6�����c*5�4	�R7'�����F��wf��c�Q��p�F�pF��i�>�b�}��,w�B����4�"h��CbH��t��>�� 1o&��4�1H��F��K%�m�&��fۏ����(�e�1T�s�P�(|*�W/�m�$�nϢ��G��K�?Z���2�00�8n�6�)�x0DW�To :��z>qH���g~tsQ���Wv�+W?RN�0A)^lҟ^������_��{����7*���w�5HO�ħ�.��ߟm r2�
<�8"�E�c���ێ钸 ����X��e$~��;��gͺ�f�_9mStC�n���$��Gd]o��Yq�)0����_��h���qfcE��Ү͑6lZ�|V�j�l�=aR����B�J~YĤ��@�,j.x(�c	����z}s�G��Fy���лf����T�ݦ�@P�@���R��f��/��J��׽��<aCX>~�5��KUDn�t��$���F�%���V2!C��oKȄ\	S�f��	��* -%�=9�x��b���/�Y "];IM�U_���˭y,����v�lR���T�3���M|���2]���
�����˘,{��r߰3n��6�h
���@C�=�J��U��Z�t]mI��3"G��C���);�x�PI�PS�Va���c��g����E���5`.Qky�y�Di���̍qF��x��2ng�$��[�t����%�z�&���cR��nnD�-����V�x)EX)p۔s'@�d��csRq)��jj��ʁlkN�ׅ�����x�(rg`)����h�o��@�v����u��a(d�fL	��Wt�I��"���B��;��NP��W0��qk(Il0��}E�K�إ�ߓ*�����e��Na`=2.OC^�j��.'�񋼂�����;��TU�U/�Y�0|Q,�=
F&ue������L�e�y�@���h4��#Uh$N��Z�������T�6$��_-�Q���X�:���<�wZ|$N�B�x�W��y1��ڣ'�R�uk�Hu3���3A?]�z��S��T��$Z�*�;L?0i�$�\�֕��e�X��� }�k/E�_�[Q[�����5�k-w��rEB��.n
9�>=	3g�N�`>-���FJ��P��%�=�6�.[�g΂��¬}��eJ�4�����V�^!�x�f��p����,�Y�a���Q�cık��6�?��H/Aa
����L���!��F"�Y4����?��N'��q#�H��ev�����4C�9�\��/��Ԇ/�9��eq�F��j13_QpL׸�M�@���4�{�d�)ivr���e2�;�E�g=�	�K��h�ˬB����p���[��m���wF�8,dw�M�;h�� ]��L�Ӽ]��Y�V�am:�������g��9q�����"@�0�[�rY>���e��m6�5	ӵ (n�T��:W'�S�%w<�ڼҴ�r��V[�<ZkV�ky���G�0���H����8p˴P��=�J����!��K���Q�6��q ���cdG�1ǹ�d��aFs�5���J�x�FM�jSߦ�X�<s�j8��z9\��p��-�^
��-K�X�T-�>�.>�g2�i�B�#ou��a� '�;�l�L��\��A���Gp=�uٛw���,����W�*��F��tѤ\K�HoN�XH+�cr����h����/z��$���QU�n�P�H���:�H�e]y�>�:���SXbE1	��k���X�4��Z$� � L���M���d=�������_/JF(M��F/&v5�`�������O�����[�ú ��jk�����t@S�ä�w���ݥ(��6�p�8W��.�Wx��м�u��G�c��/�'z ʍ0`�`i�4E���B�]��r��tnm�"}H߀]��{{ �d��k'���l�+�+��VH$8z��~jY�t��Z�뵎��wF�x��dz�3�k�K��c|���t��iT�� ��?���1Vv"L�����G� 5[w������x��½PX��������n������%r�V�d�
��@A@��u^U|�wV��-�3-<J�j��HK�e��̸tk�Yy���w��!˴�Q�ʽ�6[�o֪�3�?Gud��V~�c	�9Zo6�8�7[x19����nYH��}u2|p��^Bd�˟���	��������g�ݡ6��J�b[0c�X�<�mWS?�g��Yp�N��VH:"���
Ef�Fp�<Hn��CZ��>�y_���8�I���23Zy��B��kF���b$�7�xҬ��B�v�K�h~�Sp࠷�Sf�C5 ��$9��r�o��P��ڭ�'���U6�16�W!+����#Ē6�ڏ�%���rי�E9��ïDgO�sl`�G��YZ���xV}���d���X�p�S�3��Ł�&�b��Ð�:k�Y5���w^eh���پ��H=��o'�}��&)FX����	
��;�)�M=V�M�����{��F[?�iQ�����!�w�	B��� )՜,�=�MH1'ɐ�6�6���[:�G�).��C�_x�oF�7--�!�Ӝ	U>c�3�Z^��`�@��=�s�2Km!l�<�pPP����_��2�#�=gU�a<?��Կ5A'մ�]}߲�Z���a6�L	���'�<��vӅ�2��f  �܊.h�cL�=��ð>����i�ڟY��]6	�ؾ\4�ʻ��9/@�e~ ���C�>7��eF� �-0 ҬաB}=R�>���̵��4 ��I�I��|�)��	����+`���$XB�#�y{1=��&����{el��e֢v�>:{��՛����G����6�|���O|ڰ��gI����}M�jJ��e,uĶ��:�����;ׇ?�w����v�d{g����͙�����IN�� sc��e�|������_��#�r�Ǫ��`���p80$��X�۩F�QtPM�xγ��<�{䙬0����O�(��0�c�l��-�����f-GM�!�4T���n��
4��2�\`W�Ლ��z���'��S��t�9h{u��j�U'������k\?�##1-8�3�ن�4-��ul�3h@��͊
���ȶS�4��1�?pDJ�h嘊��׮�?琯r$hABB؇�W�`��h`2`@��ʴh�Μ�>iGxm�HT<$b�#�N��F�8~,�G�h����8KW'�ƃ�ȸ/P����X�b�A�=�Tk�Pm=��N���bn�tf��	�HGȻ���ܻ��4$zdU���u�v�-���;��U�I��Ю|�Z�3�u+����Cs�n��V5��=��� ������WIC������omF�"�ɬf�x�1+kZ>:�]@��K)�j^�Flj��G�-Fg�S���t����� ���@�(�A ��X��!e���ڹ���x�7�l���w�qhG��U��+�Y'���W��1-�C��]t��������D*8P���]l�E-b�R�海���;d{I��A��AnݿhK6*�&������gg���uů����֓V{��Y�[���sv��R~EO�=�Ŕ��T#[�F��T�N?��F�k�kJf�=�У?jY����R��U�ܾI{�:Q�u�cZ���A}:kD\c?��?!���y�m�{�@\�;n����1={���9��6!<�E�BSU�t+9���@P�:�ӆ��1*��1_=	;���Y��lZ�!j�i'���pX&�W��vsD�m�US� �V�Q|)��Bsm�.��@���g�%���f�9�7O���+py�t>�_������|y�ܒf-k"�PY(S�&�-���D�r0�T�/��1�'X������P��˧
��������mP�%Fa0����9�U����c�w�ܸ2��p��2��T[�W�I�A(/;�_Q���6̥94���V�$}3��@�S��CiۘN��� �!1�ԠRl��:�<΂����c!��9��#U��_,�#QI_ߵ��yÈ�w�xPG���,��lR���f�1���=3�7��| �q�����5�N-J��!ӽZ��L��]8�����a�}޼���6�ǘ�6�x��
#U�?��h���dAaJ��w�W`[��j�ff~�x�_A:��M�0�"�e>}{�W|*�����G��iL� �% ���T��V֠��D09�F�1'ˑ�,c��<����m��٢+[?I��8��ŬV���=�A]K�x�{<��(�g�t��.��ʬ��7��=�M.�I�(�+v��೨���l��A� �(�� .���6�;H1?&�yJ�V�����eVw�Ӓ���կ9����l�!鑵���z\���6,W�q��/�y�m��d��!�|U�	����R�z��	8J.:Q�����S�VZ^X���⦒���[s����ߙa���SJ �Q��]*L��SC�4���}���Ф��V�r�+,�*˫7:���"|� �K�Ə��G>ӳ�Gլ��]t�5�T�'��a�Q��M�WǍ<�9=_I��x��1f�^�
k������n��)�?'���ir�(Cħ�r;����;�Z+%�ͤ�,������A�@��E4"�_�A��?u�g��K�B�O��@����ib��{�F�1o��xd ��2�
�~� �~�{�0����d����������k��7�Ȗp���i�(��Vҽ5�ұ�aP-��q�vt��f�߶���(���M����A��N� ��C���)�=-+|'�Wg�m����rM�S�-i�֩�'��7���oB鄀>����*�{��]ᒻ�'N�;�C�6fg�����B�B�s�B������d�!�����L��4�8O���p����O�����@p�F4��1Z��.�ޏM�-+��!=/,)�����Z7����&ڗC��B�<�t��u�YY�������ț�16SB��߼�����(Oz,vΠ�U]g�H���d�2���?:�1s�����K'���SI:ANj|��+sA���m��Xػm� �0�!��0�C/�2q�)֜̎aK�9������?K|�����O|#�@C���u=B=�{sY�~*^��n�ԁ�z��ى�z�0G���ZNo�h+��Ѡs�u���K��_=T���7�9";���a�$:ڙ�t0h}*9CW��=��x��$���^��Sm`���}���Oè�*>����ע$�rA��yn�W�ƍ�r�*�(�YFr!�-Q_��E�AUuԱ��f�';p�C�BR_�lx�-��"D1� �����w*݋�_�Uc�g���!��_>6&�X���М+���LR�d�zQ ��F���v9HK��1�o���DT,�e� x�VOٿ!a3ʱ{@���
�hT�!_�Ʌ�Ǿ��5� eNy�6/
�j Q��J��P1m,��C���F�:��B��(����Zv��"�]J	x
�p�e�Ԋ�
�����d�"�`��}�>��6ꀃ�3?�I�f~���)��B�W
�{�i����W2�_�)��*~jP8d~Nj��g��jT��j��!�	I3���7�/%{�Il��yWW��s\ ���խw�Wa�����v��y4���~�B����7ב&ɡO[��O-n����.���i��e�Z���Q��a~,G�#�n���.)�Յ?%~W�RH}�����ƪ��2�x�=W��-� I8�^5�#��t�Έ���{���j���F2�x��vϮ�J���͠C�n�T;��D��A٩��ǣ�|�Y���ϼ懊�w�9�����G+��a#�P�8X-�-J�*̗~1_U�aĈ'��H��9�#!<|�{DO�o�o�om�R��������=Rl�O���CӨ�ܤ[ca ���Ǆ :"���/�9S�B�D������yc��V�G�u�b������lq��=��EP�Z8�������X�V[��s���P%��f�w	�[S�m�(I��i�j�U(>4w�ЀV���I��؈m�XK`���X�ȕ)��'g�G�p�U7����IT�������>���JYJ���XߩC�~�fԉ��+�	#����ֱG�pb�Xi���L�Z 7�PK�%&���x��o�(ٍ�����^�9��cd�dO�z�?W���6����bI���#V\�A���2�&t���Mޓٮ��{: ,T�{�ۮ產!0�c�	&Ii��K���;"[��_����˂W�Mu�͈�Bd��а��hU�ͧ[�7�� �{�g݂����\e|�S�~ל�HY�*���e���XM_.�~Q�	��d`X�
*�*�L(�5�)��n�����T������"7#�؈On6Kޑ/�=��3~5��ܔ��'٨��j�rW�3&��@�G*�.��5�[�@��֏}��\T����#ۣ��]�&�⏿܌��5�0�]me��B8��9��=��6r���o�6~�^�z�J��y��`{HO��J�8����됃��&8\\��.�Z�F�;�ܥG0=0_��~�*�^�xc)�1>�iGT��R��غ�^��n�k��������2��L�2�7�N8��i���2mg���q��,v��S���V]Tqd���f嗣X�p�({��4JУ|,�h$+�J�ꩯ��b@�Ok��<�L�����:Ԙ��71Su2���J����U��z��5Ƅ�1An����KI��(y��2�P�� �ƒ�z�QVϩ�����@���z��"�E3�f���a=��CÛA?V�	��*���-��P��뿠�Oih�ai���s�ҩ�ds��V��R}�@J?u�5�����;>�aib=���{���c�&5�1�>_�݅+�ԡ��?��p�(�x�LY|�u��ڧ�a�à�|�[0J�+ZBtQ7�v��?�t|��IV��o��Kb��b�u<g]�5"	^���wy���G�K�w}$t���Ӊ\�Ec1*�}c�6�! ֲ�9N2U� &�.g��f���������� ��O������ﵬ�7��7�<�9�����Qs�O�����dz�]�h�a-�<{�㿷����v$T�F�h< L(���,RVz0.��pe���[V�Y�I�&�N�I��)eIa��A�@}�j�A�����v �h�2�W��_�F�C��j�$!����}�D?�\4���4��U`E]7����E�\��W�F�6�&1��Y�+K�n��B0���0�	�2�S�S��a��	E���G?͕�C	Ⲹ�aa����N�q��]tT�>'�@�l��]�R���w�f���BG(7�"�*�*b�1������%(�4O7o�t�2������F�LA,�^�t����g#A¢:v{�χ?r�M�$��!���n���If���a�gC��;��!��Ar_�i3M�������&��m�եF�'b3����//�U=�����������$�{�A�K:���LE	Hw�ڕ
+-C>x~��F���\Y�y��4ۛ�!�ڊ?��'�+b�� ?(o���tY"ϙ�A�m���L&%��߸\�t��z^�.j��B�üO���_ ��M�~��Sr~�e29r�!7(G��Pv;aYd&m�E�������z�5=�H{^n�k&�F���ߡ�.�"t-H�� `H�)�ַ�&�-�}��N�ޢ[�?��>��z1J��۰^	��U�k�x�ǡf���0�s���[f�rh�8q7�����j�Sc�!L��GO�I+�>��B��6a!�/�L{s;%(/������<G
����c�@V̎�i�,�Z�r˪��?�u*��LC�j8��5��E���ϕ>k
)�Dg.6!ש 8�C���F�a�#�!NJ^�橐'�z)^���eNFOK!.���Z��9iղP����ֿĤ�6�V�rEd�Q����tv��/C�e-��𹹎m�hr��"~�V�������B���K7�����< =;[���>�.�=��\P����P�fҜ��^��o ��N,D5{�>�HZ꫏RvJ/��8�,*�����JB�ȼ?�;���)g��m!�P�:�	"��eM�1�"�Hgq�q�?]�	H&��FC��o���č��p7Mo�jvwB5M�֍1�b������-!��0�b��\x>������[��*�z��oT��+�׵�, Ü؝]���v��La�2���3mͩ3��o�������GCbl� 2����:ƦY���0�������g������}���n��	��h�&��-�#�A�e��q?���{�~wۋ��{}7����,��� a�$���kI��B�$��E��&CN/x<��Z�+��Ծl5y�{���\*^�c�rQ�rw�+��q|�+��!����z��w��C����I�#�t�]*�6���9]w�������C��6�?B��:I��k:Y^����dCW�,i3+^�
ۻ@%������?H�}���ںk�pxB�?<��� s�F��D-m��L_��?`���D2��4'J`;��o�w}��|q��j��.�C�8�E��/ka��vB|�9j�����mX�f���Ae��z�wۼ����15R�H;�]ܾPG�AN��i��PNkx��8i��Ǆ �J�w�@ڦ��%K�67Z�����l�Z�q,��n�1�Q�̐)�W��K�52��d���_|���9����+��%������*�?��s�H���it|Qv�J�i�9���]e�����o��.o�K0<3���S�����d���2i{��dow�ӓe*+vy�A�d�x�i{�l1ͅ�s
3�X��*�l3N8���X��(e���9����E�b8˽��{�O�&tѤ�s엪4
Q�CU�Y!���Qp�`B�V�=�س,�G|�� �#݌�&�T�������t��@݌X��膔��Ԑ�Ͳ-W�̇	��C���2F�>��ZN츥�C�?��ڊ�s���A�C�tr4�̝qc�  0P�e�CFz��G"�
Z�i��0x�$�gW��Of�q+ʂ��� �I)`1�YܕB̲Z�h��^̽w�ə��Լ�},І�,;��1oc��ߑ�1\$k����[<�	��gm�=5Y;� ^�"e&��W��/��@:d,���zJu�w�0諃������3���uu�H�(ı�.=�_��TX�Q廱���aXNU/c�Ie;52X��A��"{n���ZQ�ƻ��������s�,��$^�@$jJ��ka/�6�xl�0<l���Qk������k�m��us��fu�Li��#x���뛂-�g~�f^N
��efl�"3��@p�Q�Z|F��0Q�C�����zap�@�E�Sk��mcfZ��o��.'��{�0��f�`�I��EV�v��]�oS����� 7�3ޮIWkn	�J�Pւ�)�I_)��qv���.���`S�@��4��Z�&���� lh"�u]Ļn8��a
��L�x.��˩ oK���a6�|-d�f�֋v�_~�S�̚�)ڵ]I� ��_����N;#0�����V�^��@�g1��R~�y�5.m�<��DM���=I �S*����f%DE8dk���-"�� 
��9̺%,� �7�� p���u�ã9������"�[�Z) N�����
<�W#-U��μE�i�,���z�搿�嗊�GLr����r�|��je���[>�^�I����0.�v�GQM�od��13�-`��h���lw��{u��������"��c��G��yY�L,���H�� x	E׿�}��a�M�]S����T�c��YȐvj�XЩh4��c�tuʡ���}����y0�����h�����X���s�tg��I���QE1�B��,����
ӱ^��x�n�,�Vh�@%d�
�Ggc�a {�UdM2O�h+J�o����K������E�O��.h�NE�b�T��ɹ�.�
i�'K�K���GJ�%����<��Gl/#�����Z�Q`�����?g�������&\�xN����?,+�&h{�ْǀ��ۏGYE���}��ꂼ;�/�0�ƆE8��o��-�X�N�>����]�R۬<bv9|j�*���oR�2D��lqtZk
�������Ah�(��JK`�����J�[O����
���*�����/��د
��'�⺑Z��ȝ�{(��㱔������V2m���laǚ���W���?Tp�)N}iXA�!M�͚T�ׯ+|
�S�u�&�s����2K��2k/{+?0�dkx���-�n�(��n^.������~�[Ѩ�;-���T?�'�K��+�t�y�.s)��]*&� Fs0{P8��i[N��_���g�h�@@J+�4 e������aZ����u��R����v�2uB^:�|DC�|�����iJ}��O�q4�,�&�]��������9Fa�`@��;�]�m��'8Gؾw*OM�x0>�W���V�J�����*ק�U3���Pl:��!�x�y���(��A�J)��(�2G�ԥ
T�̬���?F�&�Ww��3��7[�II^��Pz�!��ɇ��8��6D��.ʴLQ���+.+��x�c�)d��_Q� �ȍ<��-1 �~��2�`�}["'�9��<�	�[\�E��T�.��3�9k�i{���!��cY_���W����֊~�ANg��f�Tೣ�T�6J��̫MUn����|�1sml�{͒�4>?@���6���&���d%j��R% �R���Ż�J,x�L�>�J;%�4
���JZv�Q}$ �y��N�G�sޣ0��uU���S����F/���T3��dQ��,@�JȆ����"����B��y��l���2�8ȄV��F.@)ߍ���}��X]{&��y r�73˘�f�1W&Oo-�/���X�x
3q̢EI~�t�+ݣҒ�T�&�g�"T����d�����f�t�8>ϑ^%1Q�H"��:?�o�~o_��\����������"Q�.](Y/n�o�U�+������/��Rp��.�)�:��MC�����p�P��@�6�#��98x(so���5�5@�	���9���}��q�Y��{6���^�4��R��ΞL�u�a!�
�]5rT� ��R�{h�BF$�μ&^���K��, ���C�"���7{
T����3�yh������$�L:ߒ�3��v-���x�:�U+6�Yɴ�v(i��R�ofQGO7C���Qs���K̟	7ݶk�-�%%��r�w�18�v}��4�6�f�i��'�z0��b�XM�����,U	��zu%oDA���+�[�TE�%)g�'cZdE�R)�r^9�b�����g�H�0̛�������|�`��V6��4kN	&]���h�����;�|�(�Ӑ,�x��< �^QYe<��n&�#W��L����h�/�ŵ����u`֬�u^1�8u���w�aE''�ax�4�>.�f�{�n���0�.��h�~9�)q�%�no���dG�������=Ơ��.�N������G�����>)@y����革q���pU�[n:[��r�#c�@�i8�	���5m�ƃ�{��;��>c�lOq�P��O)�$R��1����|5�/��
OA��sDBj��x�uώ`�m���@����i����v��l7V���XHLS�~�][D�C��ddHE��������GG1Y��\2.o��1h�Ii�p��/�)�G����|=��a|���I�r?�,)L����H��`��=d�$H�'�ӌ�}����9/�X���
�mK�!V#d.��k��]a� D�|XxI�$��x�s���/��Ro�����4���Rݾ~�oF*p�L�B��&�=��ms -9�e
B�;�����~�,X�U;��������w-���~�������Μ*�ݶ��˦�7:y��*v9�ΊiVr���^�5Ɂu�j%쩋�HY�dE�Jjp5���3����Ú��~6��'���h�V� Я~�_6o�����mz0��'|�ɖ�P�oN�l�M����!�v�V� _�#@u��܈'�GAy�,Zo��a�2LyV\�'/��j��m��\�T,��p���u?�;(J���)?nJ�N�c�L�3�dA��y�R��&�]��'Z��(�q��)n��$x ����i��0��C
�!�D�+xWu�P^8�+�'K㲹>�	e8�BI/(��J�ι��)u��[��W�Ӝ����h�����Sj�8wt
B�SAe��@�����:��'Qc=�vz�%��Ue��G.�4%g��O<>_�ӗM�BR��'+6�Ά
l@�A��ƫO^c_<�/3��OD\ s��L-L}���R�~�R��Z�k_�ߺF B��������*E��ۍ���V�%xiz#+0�x�+��J�Ml�-(dHG�4���i�-ܿ�$�
O�:e�Y�I)9����7�v�uIW�k�J�L�peY�@�\�Gzy�t��$!y�T�����<�;��x���%����U�ny��94���ߋ,��4G����˕�8lb4��<�3�V�z�.n�����JX	�n�;��u6Ҋ�D��n�����dd�}����C��BQ�4��=OZ�Rب�_c|�fU����r�r�(��̦�|��>���R6�	[�1�����^1�<�Ȭ����V˻ٱL����T]yM�Ƶyu�1p%����S#�a�p}�5��1��u���EJy�=�����R�p�f��^��]���.��WJ����#��)���h�3̙AK�l<�toVeOK,R(7b$+W(}N�wg�ݾ�8���E�4(|E��\.gH+3#
_;��D��y;���V g_a�8�B~B�N!�)�=X�%=����@i�N>MZ�������j��X����x���������=^�X�����Mo�Jk�riE!�<�PDU8�nҜ\��z:�@�q����O�X]�Vq��ο/Ҩ+1��D�I�e��U������K
�Ν����Z\.�!��G�����x]��j#�jZ7��wO���+��">50dR�w2'(��r�EATw�{��.I�N����H�*��� �&�¨�)a�X�pEGx<�q����V�]���a��m�h�"�.7X[c%u�Ï<M:��5� 2�R+��B ��9�kq��n����]��E�rS&�1����t�
�q�}qq�Ә�2��3�"B������Q��u���c)^A��ֈ>�3ex��-�=�0����<I�h�·����ٛ'T�z�6�֟"a �>�]������=�G�^�r.�C�cيU3�a��OV�p��,iđ73�G}=��St=cP�(Ĺ�8���Cԏ���gv�w;������IxI3H7=!���JB˄r8~=w��Ohi)��ƓbT��/���I�e���;�����.#�����o�'���o(Gi�P7�O��e�Dq(i+ ټ@0x���}��>i�����Gk����Z�>B��i�� ɶQ��s�ׁ���D���QUuU'
�c��[U�5�&j�m,*-Rzr�6x_�������SR��-��I"'�Lf��owO�q�tS�=Hs�n��s����u�+�?
?'eB�W�t޲J��K@G}
1��p����Y$;��P(.���0_�hg��	>�y�[���A��~�ψ���[\|�W��]�+�k�5�K,G�/k
��rD,��������Pe�U�d2l�:ؠ@�#��-ً��EŁ�ݐ�$!�����a~�i�Zc�w�e���:5-g���s�����S��-�?r҄�'��d�o����jM��'�>�?y�/~��=�����j�V�_�-=���x�v)	�&�Pi�u�*���`XF��ID�`Gm-S�9ރ���u��Q*���e#Rc0Q�걌Gg�{��4V������$Ґ��n�"R��[�[�ꜥ�p�,����wznD=1e=��c���Ƅ�rN�}��!��!�&}0�	*�ϳ��Ui��
"�(��lH�{9�k�~���d=N־U��kn�tg)�Y)5�ț�4z����Ԭr˭���'M�Sk�>�w�"�)���U��VHUw+��,����^ͭ<����i��$O��R�3k��o�s��4>��˚�/�����&+��C�^wf�95gs-��w��;��	�]pl�{�MJ���u�a��P��]�L0�ޡ�һ�)��&�'��K��VX�V�&o�x�C\�՞O����Z=O&��?�h���tn!��-M�������.�Wuzb�+��GEXΩ9w���җ�:��n&X�VA�tC��T$R�(C��~�`�A�>��N��.��8}���\g�>4J�VB+@��
�bd�xÛFg:?]o�B���tX�- M��qn"� �o�[#��w@ue�
�	o�fZc� �j{�L�� H�s1�z����%�ۜ�B����-�TM�G�w��Di�pa�J��@��te�<!��;��}@3K{�~(�h@�$���5�wG&7m����=��8,R�WO*uy�?������U�ݭI���r�f�Y_�+f�Vd9���ǥ��J��㭄ns�_M+�������Tcg���aaYXB�N�`���������0R�(�a>�e��,p��A�P2{G�� WwiW�<��\vHLl��v����J��f|C���q�O��L�'#�;4�z�(��&���}�>	�5�����ckXB&�0�<5�7�L=�[����8�g�O�T{�A$�y���T�%VM�"��>�7���5����;��N��mp@�Ƙ/�?"�H��g5l|�량{���n�2�p>�*^K��=�a�,T�y		��z�:��t'������n%���F�Z�k�����t��ʏ��0�&�A��qO�n������~a5���q65�Y�R�	�V�gQnО?86��x�^D"9�PU"R.'N2��� ٔ��p+oB+�����O�o���
���_�eyA�ŗm���M���\�I#��?w,�D��ʍ�*IXEW���U q����牖@!H����7��Z����pǼO:�@뇂��� {�c84�љ�0�<r�Q)w1�U+^F�A����A��0p�0�c�(��cWONdm��Q�A3ɾn�T��Z}W��g�k�p��Ң���fL��ǐ�֑w�Y�L��BT�h��L]�,�|��@5m�/U�#5� kEfN�<īJ��h��by���
�`H8iq��ˎ�J+qQ#��k�m|�=��a�5��y0�D݈Z�è�A�N�jI��"�i�~�U�;�|��9���a����՚�m�Џ:k�k�J�y7?��n]�]�#n�`��-��S1���H�:�����o�0��s��|y�Cqv6Y�M�� (��CV���N��>Ҏ���B+}Rη�z�f�P&q�.���M@�Y�
z����Å�%�bPz��͑���N��a��5
b�E��̤6m�䝐i�q0\$v�_�bu"JF�H(�v>�U�np��S� �AW�?i�ڗ�kW6�2�ۜo:m(��dSN'����#�� � (�Ϟ�*�cV��!	���s�����q/csP2Xq��V�9�cYu����b|���J࣬c�`���tB��|먨�q�PfIt�6���(J��Y�7������������`�>�&#L2@g_>�=|�O�.�ʹ����}���N��ne:�~ݾ�I��&z��c�k��x�OK�f�������S�+;�~�ñ�:�X�%sS4�d�8�.��
Ջ�vn��*�_������p��>2�yNZ&�&������0�"m��a��zN}���
N�I\�BZK��xp��;GZfhy�:͓���p-6��riN%��{F �Υ��� @_�W��<��tQ�8��
��GH]'�l=|ؤE�X�ه�Ҧ�Tn�D.MP�u��wqWz�oڸ��9l:�x!u��:�S�gX�.`��W~��"���u+�.C
�/`�0�6�QÙ�}��j��j;�S����穧�Y�y�5�[���pF�u�=���A�R�p&8�R%��������l��Xߟ&"ӆz[w�Æ)��^��%�֓ɟ�g�Q�rg�����	h	���`
���P���+�?1�2�-�F��4�cY��[�F�w͍7*$~���a��;��>}Cۉ���o��?K(Q��Z�C�������o�FV=Q�f�77p+m�Gབ��41���y-x���_9FG~��̯>y�Z����*$I��L�H���[�ܽ!�{���/�Є�l,��<������?j��cOFG�S���"����g�`�8O�	J�~�z�Y�A����:%O,��mQ�	K	̀C�㦗1��|c߁�8?ՠ��u�|�)I�!]�rח��7k���2�XTݙ)#��1�EA��!@V���*	�;{ƻ�� �cM�>�,�L�zo&����I%3�M���&�Xj]�9�ຣN φ�� yq��8��<�"�f��Q\���͘�<+�@�" o�O3X�=���.��mH	�Z~�"��saUT�'���c�ܓl�NJ ӂ$��{�(
�_ ���p�y�BmU'?�zDX&q�+r�0�z�"3�Q����w�,f~Fg�H�����ƀ;�=��sM��NB3y_�*� VȢG�u*)����"�mF���(U�_*������$ȏԏ��U�'M���G��p~[�1B��9��[�z��(��^�N���&2��/��;Y��O��!n��V�K�<�����7�.��4}uٔ|G�QS���#�:��}&����J����{ m�6X�|3��A>���!��4�k��Yɧt ��N�'�<�Ʃ��-Sb3��x�&i>�q ��.>d�iI���TRf}��[�d��3�tR"BO���s6�M���=�8�ˍG�����s�1S�S�Sc�@t��p�Ma��{�ŋE��$�n����$����{���dLj�=pY@!�w�i('f5궪R��¶rz�EWZx׏�����(��V�d-�ޠ��O7�_{S�|`t-�%�|B���$���<���=�'z���a~Ţyd�eۇ�	��p2)l�~��:��s�m���;��ԑ,x&	�:����{&¤ɾ���
�B9e��y�C��ܵ����#�7��4U�>�n2cKdMR���V�.r܋�+[�Q�>�׭[�,
���I��R��paR�LʁN�.�P�?����=�f�V���f��(4�x?GW��J�H&#ju$�I��[�r��Ֆ�_o���ܨ��ͷfb{~���J3���gZ�=�y��#)a,9��ώ�]��.K�V�*@߳5�D���j��d�`�'&�ð���In'���C)2��9^�ġ������/vde;�
�QI���׌!L�E��1ؕ��sS�!5�LS������Ճ�Q��A�(��JW��9��Ha�n-i@Q�{.`���-��퓘nMK̵���OI"~L���R�l��s�_�{�p)�A�:a�B��K'<'c��'�L}����o��Q&��N�)@��8��.b`@M1�䉵�CB��~��<�U�{�VYU���U��q�]��7U�`���a.�몏pO?���C:�u�)~:���m���%���x�S��EH'v�y���
���@򍿒��N�n�uE7$�>���Q��Y� ���8"Hd�0�	�KY̘�"d�1+�\¾���<�S$�Y�&�L����X3�UԈ �ϟ��iGJ�Ќ!)#�Dv �>�����S�_%�`�8�ڀ_���Y8�% u��Ϣ�Q�_lOQ�Q�Z4�|�r.WtM�7C@��#�2q\hކH9v]�� �(+���,��99C�[B�򍴃v���[�Y�L?+��j��7��"w�f����Tc(s[���LV����C���n��=A���s0e��i��0ϋ1>�,_Tivw�o
�>�+�Y�J�	�auj� )��@XY������5��s7}�$ c�Q�E��y�� B~�׆�F!u��r�!���f�墇F)@�L��Qr�I�7��K�>3M=U���R��|� ��Rv��~�۲��̕���PU�'�u�V������s�Ho���`m  z����q	�?G�?�nM!��o�)w+�n�4\�R�����N2A�_AdD<fd8��R(�����{�ώ �B�hu�Ɣ'��p�w��h���`�.>?�m�s����$v���]�S��W푘�(z����n�'��<�ɝ'�gݫ=L|�xɃ\^
ܗQQ�9wJU֋�]e�S�wm���~�=�����z!Nhs�D��Qg?I��g��tI�xv���녾��z���B�Y��Ka`n�#�M��S�uZ��9(����S�����uXJ_�mЏ��Bg�/��u�+r�Y�rH"�����d�=� ��t7������zv2��&B�6|ʐx?� ��_e���;���t��ؾ���$=j�t��r�`M�<m!�i�sa�G��i��8X�L����+n�19ݥ�	���ʿ��8v�Q�J�J���h4r(ed��W��f�Y
�|O�ʷ:J � �^EyL_�|�y���e�im��e.�W�U���T�F<t(���Ѓ�M��f�;��>d�C�J�j�5�ZW�jBI�ְ� �54�C�l>>��5V�2~�4��M�oUf+���,��YX�:7�v�l�;�ͨ�B{ŋ��63�|��'���=�J!!9�I�7�F'������&�űP���_̜���D�?��H�P�<. ��>�G���F%P_47H���@]�AH�xE�!%������@�m�-�o!�$`���m3�*��~�M�5�j�O��T��3�̪���h	�ot}��?�1/��6p��٪]��צ֦�;o�u�X6��� pV	���j�����D����AF��$?��K|�x��ua��vN&���Kձ���E�w�qcR���U©n] �
�#7��3�㕵��V�jD�;�w�r�"�JnW��+SZ4��<�yy�)PoTnK��t�+�!z�ڷ�9u�z�ᵐ�R1���ؙ�a𼊞�����H�u�6N�؍�,WzЙ�t�Wa/���s_���o�%��(�Z�Vޚ2��Ԥ�04��Ҩ]�?�d׭\��nk�����n�}ܤ��l~��>j�d�5��C�8M�z��{[I�S�6�j��� `�d���ik4�8�:��è/v�L�8?�M��7�p����)�½�?��K�ܥJ`��V�2)�dD��:�P;�s�/W#� �I;e���8ǋSQ���}�o�AIT�Kؤ���Z����b�i+3�qn���̬T5;��i����PKxm 11��v�f��X��{�W]p������5>u��a����5K�*��nsb��8@���?.����LZ����|����<����X��p�#n��A3��F�Z�_6���XM��c�榦��[�U�C�i��y���ދ�DA�|�P��L�p��9�޹�V� !�#���Jݑ `�X�%\������Cw�J'7l�&��q����ۡ�?BÁ�W�hmV�
�b�yf}��?�Go���I��5l�l���^��^s3��������(k�hW�_�`=f��*Ͻ�3�&�ͳ3����f'�PG�L.�M��z��|X�4l�<�#� �Gu�C�
E]�V$���oO��`��%q7�Pb܁&+�Ť1�"nI����B���4�諬k�^y���Z{�����`/�,��%B�\I�a��\R����d�ҡ����_m4J���,Omp�%�������Gu����36Ԏ�H	 �=O���g\dht�V���O����
θ.��څ?��`�@����K�:ͦ�}���Pt>����Oi�Ss��5$Z�Fֶ`���Q{�\aeo5S�v�]o��"(�!���z��׆c1�&4���+ґ-JRu؇Tq��.B��ł������]�l��G^��g�K(�9�����ğ��I/�5]˺ݞ+���+~|w{�.���V/P
GS)Y)��sڧ��j�P"'5T�1�x�փc��Aˀ� �uR�������(+��x�ut��}<���`Uw�*d��֊�k2�	:����c����I��)/�{����n��SI�֚�Rj���R#����E�u�E,�����r���Q:�፰X)�����V��,ZU�s8,�0L!h��DVҵX�ٜ�9��QK낂.�������6'^1��-S�<�K�Wu���#4sY����V5Yb�h���5���>&}�*�f���>Jk䕹-�{$�g���|_��붬�k�(!�)Q�^�B�'Rϟ�]ɓ~�*�dv?A�wo�sU��c�jBtŴ���̝+���4
�o�cP�V+���<�����[���$��]�&^�sH��+HT�BZ�����Ưj'���ʶO"7BwB?�2�r]Ry�B�Gn���ܤ�O��i�O�(d�ǖ����@#�ߦ[W�y
������Zl쒉�i�K-��V飖f�fV��˦V��{"�̼O�G�J�#BwN{D����׍	��sS�#%b�&q~jl�ԛ�:�_��,O^�����^��eM嘯�����D�x]�T�4�>]�=�~N�9$���S ��W&󌻍�V�3r�[�^�?ý���q���(��Y.e_tm�`>�J�602EЍ3@E��T�Cq�;����O�? Pg�5�s$���T�Y�(��1�LO�w��ֵ�%@{�
�t�}��:���a�~e��K�T�[�ɜ��)�ӭ�X�z�>6�2=$Wd���+�2Dt%߶M�WɩnF��甫XkH�b�)�<B\�`U�@�`*��{�`���8�ί{^.�����o�
���?y%�pӢ�a�A��o˹�MJ��F�Uh�ì�n�b�+�v�SjH�8��\wf�0J��$�a�{��%u���hA����*p)p�E� �J"�uJ{(A�u�ڙė��`t$�|;��h~�7S��!Z�Y��ؔA6}X��:�^hQR�� ��W��沊��Z�i��جK��X3�d�ÿS
��
�w����P1��� � ��@�;5(#�_���������������v{ŝcBi��~��������e`�
��w�U�c�l��]��C�q�� Jg�rQ���#�3�!�{�f7�}��h9�ԩ����~	Ly�T
�zM1V]~�Q5?�� u�#ze����$�CSހI=�l�j���F�t�so�n�<08��i�%��u��=�Uz��9���G�׌<��8KE7�VoD^��'�Qk�h@x?��^�,���C=����r׽��>b\bWJ裈�r8�S��YD�fLoc�D,��~���<}�ܧ��k�f5�;���;�T�����7R�}�D E[�Ɓ
�փ20h
�Тvλ�{[�c�����S�ۊV�S������)�)�\ ��{�g���e/x�d�8�g^6�9`NP����L>R���*X���ƦG�5	A�c���
�B�4�S������~�2L&1�����t9�|&��r�O�:ۍ�+��F���WB)�4�9,�E�z̈́Q�(��j���� ��)� K{y�
qѯ�\�P�%@�4��ͣ�	��˕G#�I)K���m��S憚�bz����d���Sz���U�M��Ȭ��>#��^�� ō���7���tY��,��xth��si�O�dz>uC+l�.ݩ�4V��O�g��E���s�B����@J���<�-M.;�^t	����U�#�=x3a��Z���/���{$�%��5{�`x��ѥǄ4�[k����n��w>b�,³�#�d1��_��1(׃��Co�!COD��
@���7�.�Y����Y�T(3�c]1C*�Ȓ�������f�pxx��s��������7��V�ѽ%7Uݴ�i�(�;�40-2���Љ����h�uӥm���\W�4�p��Qm�P�\^��E��������8ul�i
+�����y�X7��Xn����w��b������@��L��X7�(D��~]�+8�3a
C��¢��.�;w0S�р��8����z/K�,��.�ȊN�{�!V=L�`Ë��<U>y��"C2�o�JsZԀ���]?�S�(�Ԥ��*q�C��oJ�: ,R7=�j	����2�$sw~Sb���ͳAʦ�����8��{����&
G���P��&X�`�+�ֈ��x��3�����Ny%�y$B���N�<s��Go�4~]]�)�D }����������yi)߯,n��@=_�)�Ml!{8�X-�����m:9�����v��Φm�c.�����fp���B|�����6k�M?�i�J�X��(6�rE���ȓAL7jo.��<�f���L�.B_�(���������9;Ay�{2F��V�����hK!I&�(Q9�����!	�`ll;��+2�^L={�j8��=Ӧ0�������V�K ~����(��O�j#ߥa��ゆ9N���h��s��f�3��(�\l:�olP΁͍�$rE��:�"���B��vfH�ѳt�:\��t.���Uz�������kt]�hB��GE��%qk
���%�U�ΔR���Q`0�2:<9k�����|�28��ZJ��O�q�ŉ���腻ڢ
��a�����UԄ�E�ǈ�G��
U�w���8o���p��b��T����:�.��0f��_sq�)j�1\kh
��i:}���9�ZsHz��)��qvS�xM�%2r����5aw�w[��6�C)�-�I4��w|d2b�"����0�����Xܬ���G'KA�q�~��j�3���pX+,�v-t]\k�!G�Pf��p�,�u@gEu2��?��n�I�l�C8O���e���CL�[)r�8Dt^X�<��p$�]��jk3� ��3�wņlj�_�O�І�\�2]�x*B�C����<��mP���s�f��A��k�*���:�q/"�?��S"�*1f�����Q��7�چV��@��lD��	pơ�ߚ�{������|Ŗ;T�/p/9v�Ɉ�ɤ��q�z�3�j�����i��&g��z�R/� y� ��+���.E���}���G\���:���f�Ι���JO��a���Hƌw6���|���|����>]��.ؔx|�dRc@%�n<�����=���$�x�=h,J�z�	�3��|M�IE#�2�U��Z6�B[⠳�Fk`�B�|ú�%>u�S�"1�P�Ky޺�ˡ6��!��m�J"�>��U��ۄ����#c�@�&��t��J��^�����������e�g��n�(�_���l8?,�UX`~:��Zy�
���֮���l���DP�L%e�d�Q��d��P�p�������'E�Z��0d_S��_��W/�k���D�`�'���{`��U�H��J_k���ZI�����#4s\;�0�qY������� d8l����>(��E�
��kV��@����~к>��}��W��M�7q^`$���� f���G� ��2��,��=)��b�����C6��ÃA}y�4��:H�U�>��w\��ꛘ�'%ăĘZ�9���p��m?w*s��ӣǝ�� B��F���J�)t�_'2������r��Uy�}�a�x�:�b?"����)���L<w}�1�q��}��@t5��^|-\��h2���t�8mpsnS�$����/������$�"9Ds�E>��ެn��^s-�J�#�����]�� `�wvtt���=���ҵ�y)�� CV)��,��nLhpI�JAɤ��R�vn�h����J�Ν@��pR:�\����+����~C�>�<�\/왩9��M���$P���l�@��p�D`.i`�qNK�3x��n��[�D�5��9ZQ�OX���p.�䲈�@ȇ�+]������l�O,������i��e�Y���@�53�\4�6��ed�e���賅i���V�)��X8���1-���$ qbsŜ0��'d<͈�[�^�;)��2���}b��yi�O �y�m�{�n�r˧���
������##���R����^q4����3<��m�G��'���"'RQRTXW
#"ZWؿ�9���� *��#��<��g�G�Bﬆ9�:ߨ���x��0�� rvMj���W (܍7H��K�$y��vkw-�?ѵ8f�F�Hꊔ�<��ѥ��}@aO�A�����hZ�[�L�Xt.�q}0z�Ҹ���[6Q�p��I���aP.3.35?)�nk�k�@o�m�5�H}���ܒe�a��Us�Ȫ��7X�a��k_�6��@f�j ιZ�<zY�m��R[,�y���+q�	x5����5 �1r�Q�)F���%on�gA8)�4�\KY�)6S��}��ӑW�Q�u�\4$��ډ���r}���j^k�-$s��.��@V/�x�~��@/ )�پQ<�v|�v���|[����a�y(������S?k~[�}��{my�9@�լc-��A�߭M����-�߳�����zH�d�Y�uL�' )�'�gc��@��q5�粄EX�9��3���i͇)D�!���X��_��Ek�W��#�^�I�G8&*kͪg>��QL�K�f~r�숍�j<���	9�(*A=J��{w�o�T�A��Ad���q����zT��y�6��Ƨ*�O�/��S}��Ѵ�����h��p�/pU�~���/��O���ZRA��
���[���ܜg ��p1�J_��JRpra�����=5�:��V��>�TٕޒS��W�ztqO) ��@�1��N��k.@��i��1z9�7��aS�u�J���:�go����u��~����
�D�$��M�_�^q�S�!��.�Q@t�� 
5� �։��H����(� ?���*u��f�ޏ�E+��ky��$i]#��K�¸������[p���o��s6غ��u�N|�%�>��?<�M�|K	�xt�,Ѡ~_q�ݵ0`���P/�l"T�����w��+��R�Gib���^mz+�񦙈�5	]+m�F���x3�ӝ���������v�I�Į���0_tN�yǪA���8?������îy;ǜo�$+�`�:���aS��p���^��V,���Ew��O�l��@�/`׻g��sr@��/�/T�vO��ʤ%��n�D'\*�Sɮ�vR����9bu���F��Uw�Y�Ԯ���r�˖�z�0��	�(604^$U�Q�xp������Xb��a��%��h�mő�����V�X#�#�Ɗ��y�[��3Mw*lt_?�Qjz��b	�"��1�/��	:���Q�@�8J�H����:DQĒL�=XQ�^`�n͉�#���e��H�'�ӾZp�<�Mdnq����b�;�˂;u^�bXA���S󯥫W�j��HT,K~cUb��[�}���D(��<�.WRў&��F���q�x�i�.�Дr+�߉	fj�jf�?�����
����D�2�'�iC'E!|ȸ�� @�6�mEJe&���;J�W�D�/(�YAG7~E�;���!݌�MbRK��M��B��-�	����;?J��fI;�-j��+��o!�,F
h�����_���M�>�VP;�m�O��Ơ�/i8�Í%���A�>WG�	��6~`�1�f]�V/��?�Co1K��G82����=�?�?m��/A�BzL���@7�m����sG�ڟ �.��vǉ�o�
_���:�+T�Gq��\SCku�4�E0��,����=�e�;C�r�`���To�P'� �9<�u�&�k�������Kx�#+BrB�M2bt��0�w��ǣ�K3h�������4�\m_��#vA�rV��q��6G1i���龼�鬭�cA�+e�B���������Q�&\+eq]��z����#&�b6��K��󿛮�v|�&� ���&���B�=�,�>�ă}o�&E�鮽�֧�V}�"I�2U���y�`��ٸ�K���6f5'Fa9�!;�p��5Y�qz���Nh�z:+���"��}J�!�Of��\w	���p�P27N /`JR5�NxD���H�
j����\����T�����W��d�����!��}s�1�S%�FA	7bC)�Dܠa�[$}%(�],�f��$pm"Ɛ��X�h�-�!z�3`YF�c�\dgL�LC����e������Z�+3������O��� QΝU��Wmύ�"�3b0�\£T#�탭�����ݰ`G9��|�J�	
�/���� IRt��U��u���@FZ`6�lS�$ج�w�Nw!	K�w�;�����X��d�С�Q^��Ux����?{M��r��9��2-�e�F��`��pꆦ,-�'	*zT܏�p#��d�iw�KW�������Srr���FLJ������֛껚�luɧ.�o�%��L�^���]7������oՓmb&�m��p�O��w����Nh�&,�����dT�����x��>-S�|h��K�<	��Mm��f�k�̽�~�8	�	Z'dVL��in��E�D~���mO�*��cb�s"���D�X͔�ϸm,���D�c���L�;�=�~�uy�ȏ�,�Cw5����3�r��gd=����.'�BL<�s�LOy2�	E9[ts[�-/���'z��	�Zm �"(ۀW��)w?$��"��QV�$����H�I��q֮���р���.�
Y�I��:`�%Q����Q��ݧ�~g>�_���w�X�����g��I�+�Fvσ23��]������%��s�N�VnOO?���ӶI����l��rz}�\\���F_=B�l?'3���?���A\���֐�i�MNi�n��f�Nu����,o��>�{R�S0		����t����mU�l��2F�46�f�I��"��t A?_�Ab'�6��0㺡� 'Mb��c*c����I���B��WF�E��$^���d���6��Å*9�t:��uY�����W@}d�"��$6d.LZ��O�e����Αr �=x�Z-�tǙ4��䤇dcϿ�M&R^)K8q�� tl�-�����>�O��X\P�5�������[�0���*�$X��pzܠ7%�=7֯�sy�,�T��[ӏ�c�trZ\���-���� 8���a����Bt�<P����t!�~�8��`�}G��ˀ�Ң9��y��ft���Wƙ �ԗ�:�+��(�c|��a�?�y��6��Q����\-�g��~��$���7�TodG��X~8{֐X-~�D��?��[�z�"�
�u�zi���QN����c��S��LW=#s���I�Q�:��,���l�,O���&�Q�����>��3���X�����.�c�,h�!L�C�0K�-x���]A��6
���Y���	3:�*+h�R�$WUbJ�i:������
*$��*����N��T'u�5���:EZ]$*Qb%���W7�z��ɉ�L���
��>I��A�W �3�w|]s��ڥa�|�G؂���|[�@^�c�@�mr�� �Tl�?��hqT�S���֨��.*�~�Wj����Ђ`_+�S�-� -,�HbefH/A�`�z�O�B�ʚ��"�0�<q�^���E�� ��47��r��1��#��ک���;�w@y�`����V'��u)�$_hΏM��X�O��њR������]G���켣4I�"��+W�UxN�鯭�r7E�s��c<��y��8=��h!������ǡ²���I�����
�exJ�����3 �0�ҕ���:���㈡��.	�	���&A
����H\�@�P�v1�tu,��f�/�����Hﴮ�V]K�.��d��k�X�CU:��-�
�\��.PL���]���K��[#B���)�i�̶{B;ZM�DA�,j���I�xf�n��lަ���Ó����(�l2�$i�Uy���.����	c�o2���i�O�wC�l��0g�����\��N�꬗���
cY~>`�Cl\mn�=OA��)�c��=�b�O|���&�Q+�8A��ep�:��W���}n	��T�41���/ь�hraj�e�wj�Fs�8�4�.�ˏ0����	N��)C�zFd�E5�w��ZB�x���Md4�>���ٿa�J�6�`#o\_IP։d_9�2/�hzB�F�f��B"z(-c�y���h?Aiu(�urc�ὢ�5)#q�\hi��j�^�|�#�����i!ګ�bǽБ`��.�t$=	��E]i�/;a�q$�[U~@ɫW]`ej�!�f�ԭ���-[��_w9�d��1ij�2��w����?��&=��d�٫א�O����*�E�I?��f#�in_���#>��<wo��
8�>|�>Nʺݢ������F�M���5xh��G�W �@�7��G��_��X%w�>�XU��-�M��L�-�=X
°��l>�qE��n��vZ#e�ה���kj1�bD쟒�`�:+%f�E�����K�Dy|d��A��>��� ��y�;Qz1?���������>������m��(}��,���}ynA �@I	G�z}� '^�I�Zm)K��׈����|k�(�R:%,4�frZ�t`�p�jN�{IzJ��
&��B<�op
�a���]�L,� �>&���� ������7I��q\�#O@�[s�����P*sUI�$��?/�����ю�g<��x�Ryu>�M7_��ù��4�A�%�Kt%�Oq4xϣ�����|?��dqj� �˖�e9D_����H�zjQ��c�,����7a��(��CV���O��I��������~H��ٿ�P�z�M#h��.�]�Z�N��䯐�.��'�bhoβQW�YO��=01L�>p�э�p��<�S�4�#��H ���lRt+��b���i����	w��}���~���A�5��/��W`���@v�c�H<i�T/�A#�$ļh�V�}����6�&r�G.F������mB��*�P��,���qүͭ�i��G �(�if�����`	��݂��L���9�DF1�<�.vz��-�B��`v
��z�oFC@u��R}~��P��H�'3A0��V����2�Q�R���o-I;(�U$��t�su�<ؙ�ĩ2�V\��F��(�Ji�s�B�&��d���0�ق��iQ��7d�����D[?��n���PA�>B�bS�!�Ps^h1Ҍ�����{l���������&=��Gy���g�)T�q~2N�[���|�L��G��Z �"]��Ŧ���o6���_�V�'�ڔ�h����6�.�
�>�h0�XXs�G��De�B�>����C&=E�x�g��%�t�����M�}��HN�`k$�s_{��K�WW��������ߦX���1�M`��)�%�)E��R�APX�Օ����/�@ )a�5ig�R��5���VɄ��x�H`w�h���idL��9�N��|��VU�j��XGl�H��[		$��>}��#nj��0p7C��oZ�F����h]p
8�c*�l;8�e):H}Q���'�0��!��J�pD��A͍�RE#N�t�;�ȕk����XK��(�������r�
�;��e!O� �[qp��tyi%=ݕK	8��^^�Ҁ����#k&�_<�7�Џl^^f>��^񹼉�(�L���K�c�cн ��#o�w�����fe�7Re@�8�WY=�G�¬_�cß��/�`]�P�&�sޱ�u�$�%	�w�J��o2�}�d����Sh�!F�`�m<��̝�U�����M����;��c�7����(�����Z���'��Z̛.-u�zn �s�k���m��R��O����n���=g�x�5��B�n�G(�[�a��X\� �@�E;x�3�_½����؎������hty_|�mtS���t���&���aE�Ӏ�G�e�ئv�vo|�OᏫc�f����QXzi�tU�����/}��l��ѿj��y�ꕤ��=�C����:�@P�'Õ�\(��D�(�s$��@}H��)��M��۳�����Y�2r�d����k_�����03:��O-���M�V���<"��쬫��q#�Jw��N�@��̡���Cvcܰ�݁�$z�^�6mu�\����80�	�qZa(k?w�y�W���¾��L9�[ƠI�T�<N�\j�$oN��m8�ɔ�J��U�깢O��d X��m�r�7y�S9:�͝ϩ2�&H��\�|�ոQ��Z6뮟�u��eb��� .�g"�+W38}b\�s�oQ0�����8#@2�U�PT��P�v�x8�WJ�FP��	�X��Xe�o�XI���5��MD�̉S�W@b'e��黎�!�4~wu��c���u��]ۮ���_�.F	W������,K�4A±|X8�5QG\�o�K��O{�vn�Q=�%������!����I��n
�׭��om�����=y�Vǻ��~�樶�}�c�-�FiN�������)u�a�O�5qWz����6k����N@�	񰭌�z�a�`j`by���I��0�3����Ƃ5��(��|���,�y�����⶜��ɑ����L�
Uhk4��*��yɘ���R<X��,�Q���\HN��o�u��ڥQ~���.^ຑRb�#'�˪��KX��f�z/u�ZAA�`O$c:��ds��	˜|�)����	��M������/����;�S��z�(�YC##��o�3$
nP#�u�Q���;BM�L������=>�g�f%W_6��2.��; ��"���W�(cP���2`OM���vn1+��b����6�|J���~��߷�x�Xms%/+�/.V�z5��ӳ!���.�� �ߎ��5ז���]��&��$��7���
�;W�� m��Su�r�*�:ͽR��H1���|�����L�߃���=��ޏa�͘Znfҋ�sAA�B= n؉�j٭	G�ro�T+��oTꋿ�į��Zs����Z(;���)Č�"�V�B��~+h�̠�� 0��DB��j�I�N~�� ��
�ӆ��(�"K�����n�au�� k�)�g��!���Q9�w6��Y�I0I���wĞ=ZTa��5�dM�A%X8��u�&Ht�l��-���[�fA�����w�t�<61�� ��&߅#Y
��o)�s��A`R��I�>�|�Y�+t� V]*%q��(�i�ki����T(�[�=���Xdr%���^	����g���l�ӳd��$�B�IbY|7{t�;���`�y�-��˺�*Z�^b1��v���Yc��P��_vک_.��h/(��8F֠���� IZ_��OH\!���5e�,1��:$�B/�A���R���@����O����;}/�*��LX��:�����0���՘;���)�n��D"B �,	����]Mm o~�-��@a��C�����.�z�/$@����'�e�uY�P�Z"$1�e��^Pa����.h?K�4|^��%�`>�Ւ���oA+˛�Š�W�Ou�����$�D��ڞ�� �0��������Y���L�-x�a<��I��[\)�
=??�>����'��u��}#g��&j<��zf��mzV���2��$�$�f�N�a�u�F�M�3�>�����������+�N:%�����]F�������q!�H6�/��h)���S�pm��r��{'�|�^M-�{�4��9x9F ��U\������i��#�t	 ����	_Xs�[�9����N]|
��r������(�M�y�(���o�/L�Ҕ�l�ԅ� �喀&����&+����M��H]&¹Dh���'2_&�����`�ҁ	��R�K�(���US4�To3�:I��]v��q^ʴ�q�@�!���ޛ!�-z��?"c0ah��W_qLς)ɛh�����)�#c}zRζL�4f��������E���~[=�������E��V�ǣ��/��E�A����$>U��a��?�QzU����Թ��Q��@B���+��KGh���ᴉ	U�(��tᡭ�WB����O�w�=5�5��2V�ƀT��"�1��$�c["��Z9��fVp����HE]�P��]���t �ջO#D�(�(r��f1�9�"-��ߋy��V�#�G����b&Hj�wX;�R�O�Jت�&yry8`%��Y��M\�)���O���Y3����8H�R�O�o�~����g����]���ͽ��he��m�v�Ґv�n,�R\�4��i*���?�t���i<m6�D��;���Mn>@Vy������-���Y��s��1�!�Y�͎�^�  ��If���^�w_tP�װw�>���xw���Kj<a�㕨��!�ʗw�b~�@)���ѵ���E'�]}r� ��'�}zt��t�(r�U�/�ٮI����vx�@L�+;����:��}�F��
w�҈����}OE�����͖�'m�hX�(��<9U	=�`�d5�˾1�cN�����:V�[o���+Uwi��e�vE���t�ϜBm�i�m,�U���������u5UBUY�əа1^:���4�(BO6�K��B%�����6�Υ���_ͣ�����?UO�׼|��s(�,5̓�E��M�O��A��[�8D����!��}���6�찣�C�a���M�wT=���gw��@'�Ժ��ѤW�]�!M��:�%�_�������v9�7Q?�ہE���wpu�6c�5T����V��^����4��HZ�� �x�N��E�*�x����4܏��|LŶ0;Kd��| �A����1O��2Z���0#��n�Gay:W�5�ZK��a_�p���C���D	 \�E�"L�0=�1:bbX���Иso�9���ǣ���,���>�F�1��Y�&��^GcM�5�*����>�|M }B�w%v������u)~��G�~�H8��Ez�\q�!��5�;(@,�Og���2��C��� ���!��C>�(�Ů�͟W��#�p���T��ߛ�rnf64_A�	�~D)/F�3��2~�n1�尽of".��},-�:T�A�H�-�$8�~��}�EO��p���&��pG�,�����W��fA��No	���C�=�b�!tC�EmS��"ߌc��e�φ�45f�>4t�t��,!P�}"���F|,"<���h]�Ƴ�����r���1@�trr`=M׮"����X
1p�\.^���v8�I�jn�/.���v���7���u�se�+���͂ŉ�7%{�hE0�S�GԀS G����\gHR���h��:�̠��l�V���Z�5V`�RH�q���Y(JOB(F�ʫrS���U����������
L?���sS�{+������;!	��_	a��kE��C7�]h�c����`��ў�,"��)aV*��-�����^��@�`W��҈ܩp�@��=c��ciȌ�q6�C�0X�CZ�F�xN��.VCz��j7=�p֑ro�	J��'C@s�0�җ|i�3G�`{�/���@XƮO ��1�
���\�ؑ���cN�	����^K<��6/���{)�2>2�"B�g�b�Y�% �Jf��!r���4�h;�ZE͛�r��62��כ�����)���w��Cvכ=���8D�zycK��������-�������Z���aB��4f�����)}+P�Dܛ�5�M8�G�rOr8|y�U�E���ve�0<�RT���B5;!����k䅞�[67G����G������s��xw5���[�/�p��V�H4��T��\�Cl����Y����4������BU緤t�թw�w��q�T�:��N� ��kT�w{��E~l+7)���3]��G!��V�;-hc�j1����|<�l���KR���тiK���t��|]���'^uXp�zEp���h��r[qqv./e�z�n`]�û��$i0yaٴ-�5�`�fj�6�ze\\�=k.��b'ˌ�
�r�aCR�e��;�������蟽�!���1�,zN�Ǟ���+������o"��3}U���������K����&I�?A3@��`�r��R�ͲH��X�ɯg��+WN�a�>j��MuKw��-��G�>���+��3�q��ݝ�y�{�83��0y�W#��ո��=s`�>Y�J�}DS��׻
-�>	{�������V\rǛ�2b�m�\;�ڴK������:�� $����T\��b���Ax�w��9��u� ���lM���ɝ�y����d����0"r#�n9����������h�e����kh*�Y9@�]/�o�xdV���6��Ryd��*��OfUx��Y�I5=��z��Q�7&U}&>��5�i�Y�;�!o�a��0Q��WV��?�e=\r��W)+�ԯ���3"���_Z���,��7�i�nv� l�p懀<�Վ�U2ևj>\D�y��z��mx��q�'Q
ܥ��:X�h�	��ĭ:§$�%����G��=#�#+4�`�9�~�,���Lh�a��w����iq��1�Vf��N֑�����_	���.ME&��4�+���|ۻ���k�3�u[��=���M��}��Ɩ�q�ߙW�Й�Egr���H�i2��l�@2�ۇ�w,�Є|�̜��T��p�MX��c��B2;Ҿ��_-�����m�u���[�� �䖞� ����[�>�1�[�u��)��K��/h�����i$�vTl�^.UhF�:�#9�J��Ny�q���5��4�gӹ�(���Li�ȩ���Ӣ�ph�����+����2�.P���?0���Ӱ�i޾���F����^��c�B���(��v�{�!��%�r������VPlP@�]�^�`���9�ij�ȑ��P҈
��vCU��B@Jx���Js�6��0�kp}�@���A�N�8�?����V��yR�w0�L؛�JTWY\L�w�˖4q��\�Q����s!$���T��������}�%�2�+���V����y�1�u�DLP���y��?2��D�S^jg!�/_(<��(��)J|1�s�� ~`>*�E�F��BL�#�߭�<�5�k��$���6���F��8|��i1`�֛I�������Dy#JAZ_�G��q��iCq[j����&*
R�J#Z]m�q���m��:�ɨo�uO�Rfֺu��۬~��d�5X6h1ۮ�$�4��w+�V(� �m}����Z�ѻ-�����(f��O}�]�����r�7�������3O��@�[���KO��n ��-�F�',��4',�I?�Z���Bw�]	�*�Pjs)���h��.�}{�'�V1莦���:�˵/�N�ԝ�G��t�3�]�k����٢lY[j�V��hL��䰵���YE5x��x/���8H0�fU��y���-l
݆n�]�ʾ�����p����껫s�c%JS,Uľ�)u
�]&A��I�����
,oN �E�vb�����Vy%D����qW�9�:�<�l�fO�<z.oTa�R�nb���� f�ci�3�q��ȯ�r>�ݜ�%�������$�?��F���n�>߫,���c�X+ݚ����{�3��j��*��Ճ���ƥM3��gS�R���:��څv�ꊇ��i
v5Z�8N:�fL�6�7�V� <�Q|�d���V�;���ТShRdQ��4M��D�bwe�w�T�r�*ٲ#��r8f
	:5�I�K�
 UU'#8��M/+�� `��3<��!f�Zm�B�MS���iӒ`��Iƞ�F�|�)6�'�8��:�_��;��47�u1�q��߸w"\eЍ:�a���gG7t��#���Sۃ�-j��/��:�g2,å�&�b��s�LN���x���WW�TUn���P��;�6E�F�Ԁ���K�\�i�F�m��HJ˛ΒVV{���KL��B���Z/�kL~�� ʆU�td�]�g�8�/]�m����P�Q��s��ZY$+{��<P��+
�w���<.�J�h���YI=N�����d��h�y�E(��>1uF
Yt�ܯ~��'
O^"|Zu��su�`���F��2�������1zԨU�p�y�ئW�-��"�y�lI�Qʙ������7�C��h#��n���-�̆�O��>� �p
�\�l&{�?����"62�K�]�Lb��Tv]OP7�`O��R��߂�\� ǡ�s��$!�"9ͧ���j�<0Q�NPs)ܷ������%�7h\�b�-�T��,Ѳ����Q�9����h��M'��Z%H��f#+�9��&��6�,|�Wf���5ǚ!������;�^�>�_O�f�~�D�4}�,p��Ul�.�^!���;�/��D�L�Y�"�IA"VE_7�ѓ�Z<<1���m�M�B������}6n1���u�Ht���cJm�M"�����J�
s�,t:�	��G������	aO$�d�9ǯ:W���'q\�3�
�嶂����0Nց~oUpZ�H�:
@��C��5��/a��jA0�e��Q'���sv���M#���������p/�Rx_XɁMK	9Ԓf�u���A	|��s�$�h��:K����X*j�By0!�1�*��م����j��:�|�+�eLh�oJ��(g_y���� �[וm��`�*���5�F���iq��|�*�6T!�i�HY%W*�QD4rg7F� �c�2�Ŀ\.���*����k���9��.8��	�W;���r�R-��Ӈ �Zi1�%�>$%��MX7�1��Goe��LqA�y�2��z{Y�4��l��Q�!�+#XˤA�5�7�Oe�W��'���~l���\��e?�L�!��bhOS��SZP8?�|�L8��T����)��?�g��5��|e���=+ƾ�bR�?K�k
12:��MU��''�8�HF�3u*B��������QX��V+��P�/��_�)��M�t��E��죚$!�TH�j-+��_�? �{�h�N��k|,��m�C�z`�IfS�Ž��5Dŏ
a�h��cs�T>k�����[�%��8��/گH�[T�H���}�V�渽��.yI��k=_�_�՛�dc���S�8���1��mýDl��nlٲS#�c�~���C>�����'<��h��5«K�ioWm�h���.]�|�}|.�:sB�Ȍ� y�����PC(	y��M�T@˙H���R�%B�'��^���_��.n���%K")C�>�m�)R<���U��k�Q	Ǖ�:s����	FC���ecٽ��	��0�b�2�x�B̆n5�D S�r��q�E����8�棤6�Gf���1o�NXZL5}s�)u�6[S�H2q�U�֫�!��ި$v�8>퉂H+̉>hzR���E%&_D�Vz���b�؞,��s
��U�A�p݅E�1Ä���^����V��͜A��5jiR�I� ��*�0*´	R-M��uNW$*�a��*�X�±æn	�ߠ@s�!`��1�}��C3�Ť?4��x�f�r�U���N&`��g�yf�mX���*6�+��+~�����F�,_��'G���YW,AS'A��a���]�[�A��D|"���3�T�Z�&���9n�;�����2&���L�lɓ1���5��Aܖp	�Q7+�oh"�� �O��E�Q�S@��+0l�Do��|�b�AE�a��EUWՃz��a�%h��I0�e������!b��Z���]����Ɲʴ�0�p�Ⱦ���Mvak�Y�42������ܕ���[���צ�"�v�<��Ɠ�Ⱥ��jm��DY�g�A�լ�*4�>tz�]��ߝ��4��<6-���/�{a��mB�&�n@�G�$kcE(G�>��(��Svls���M��W�	姧x(`s��{�(��� ����F&a ���~G�!<9�4H�wZ�yI����Qx�cC��љ������;��X$��T����T,@��(�Z&`�-D����\%n��GU�^�<�VW_)8���#p͢ ���&�W_$t�Pa�5��^1 n�Xa�Qg�����ΊsA�������Sm�Q'���+����t��#V��3��E��
x�/�i�{$�hK9=Ufh�V`�WM��;�SP#��K%��,X�u��R�a�9���c�.���ɤ�_���7��[�a�#*�����)0�=y��T7<��k���gv���=�	��GHJʁ�NJ�I���>n��˧M�����Ґ�ӬV����ކI\����c
[��3��dB�K9���ŸE�޴������{�1Ħ�ŷ����g�
����>��jȵڥ ^,�W�!�z�ݺ�������n���s�m0��0}a�ێ�\�'�yyb�����*5|���v�ǐ��0�ֲq)泩��f%n� _B�AO�p;T��Ө*-�{�Q0�i?'�: �+�rx�Ui�����b�mƼ��Tw�ݾ���=�Z����Є����($9�� ��2�͂��%��ɘ.d���i\9Ǘ�4����c�|\��=�|�L=+W$3b�����^@�ʨ�����w= ��t��q=�bW'��O�A�Wa��2����x����K�jaf���)���c	}�a�b���	y�Ow�_�:��S�!Ohř4>%ƨ����]
#G�r�7�,Qf���ŵhas��Q-�F��  ��w��ݤ�L]�b���Oi;4���ı�>�"������Ȧ��|n���.�9t׿V�Vdҿ�ɇ�/��#���ڵ�7f�~�@�V�>t�`cF9�p��0���.��;�w���HOaJb�O�Y���ȻEs.�J��1�3�H��&`�����q� S�I�^i��	�T.?=�f)ɂGh�g����1�X/�#,{��hF�RqG�8h�#�҄�/PxFq��`�����nOd[-9��%`�J���b�U����%���o\�rwS�T���Y��S��Q�L�͎+����y_f0�2I^��N�;��܌۝Y�m�m�Q�:��*j�`!L�D%�u]��|m��ߨ�m�r(�$L2��J�
��ٿK� �s`+��� 9�m�9+���굺����O�'4���	��^�R��sgBC����L�/��K`�l Q�ҡfii��f,��?�É��qu��R�ݛix��XbI}��j����=1�ʤ"�Uo�!�JsA�&i�Kiw�e�I'ZM=�qۈ���>f��N6i��{VU�vH�
�S(2团ܐ�g��lp�S�+kۣ
�6p���^��V���֑C(�B��rňA��]Zt8���A��#����n�-On4��E�;��-��S�������?��N�kiop�����,e��O�A����x�d��>�"xD�4�!�L��y�I,"���c���D4�2���s��Y�[wF�-��~n�ů�$��w�[ث��>g�cLǥb�B5y�vw��B��Ε�$�9���S"F����8��Owj�;!UJ2�_尸��-��9�[l%}�O�S�*�<�b/P,8���&���]��X��WX�Xg���_鍑�����Nƭw���?������Yq�J:�X:�~��faE�q��ߠ\r��
t��a�ku޽ATq`y��u&.�{G���r'��pHd���]��}��U���v��	DJ Ɂ���� ¶���/��e�r�f؀��/�\����{��ͤ,��N�����eQĖ�%&���b�o4F���8��O��Z6�Ҧ�W	4l��E�O�tsQ�ޘ�����������ʉ�T˶J���>�����I�����|�V<�+�I!�P�ǌ����.�y��#0ݢY�IHl���9�qH �&i�A23�&W]�c�M�w�u����>)ԃ?H�\��XH�t�������a#�&ʍ:��:�k��y2�8�[�Lw�����[<�1]z�Z���E�ǚ���udZ�c��l݃�	�)_`��y8�bF�<(��0��v�@�dT�ۺS�ñ�lF40�-d��wҀ��yV%dh�:M�Dc>/o����cN�D|o8@Z���v8=B"���z�6�|�e�"HR+N=Pq,��Pj����e���!����*ü�� ��<2�w|���Ⱦ�6�u�u;azfC]L�$���ܵ��a��:��s���b�� ���!G�2L�H�ce�������K�.ٳ���l�~g�m���IΝx|�^f]�G���}2Djq�6'�鉮�3- ��7��"/��IA���>:Э����l?�������o�KN�w�gB#1�y�ˁԆ����.4�^ K�K�?L�y;���O�b�]�>
f���]��$s��Z� �਴�&����P�ZC:��/��ظ[ �*0����gǦ�9_vB?�J��_�>Ô��Y:����P��YP���X^���D�^2A�s��y	*�S��k�hХ�Q���s@��`I"��!��KCm�
g��R��#3~@�|UFmQW����㌡��!2H��я�����-t>�9�7�_��z�n�(�x}�����(ՠ�Ij��U��{&?���3R?�Љ�fz6n�A�Ry%���P�9l��(zDg~x{�"KӟL�z�z���g@�Y���Ƴ����0o��>����>r���e�:�?@۳�����#��{�WaN^�N;:��܉(:�y��,������g&��E<���|�l4�S;n��.��=7�P�o7VkV�|[*''�F��܅k ���G��l�mYS]�W����M����\9u:ʟ9@�Δ�+N8L��'��&��.,FV��[�j�{����%��HM��pPvSd�'��5���h|���b����gĄL&��^WX�ZK�>�����<��.���HJ���Z}�ʼP�ov2��w�*O(����GIe�, �g�r x��DTA@y?zNՉK��Q�`7����V��i��jB<��7R��~��k>�!G�}i9.-��g���5���`C�|�g����V��T����]�a!Pݾ���k�y<s���њ�I'�����5�`�?2���8;��6x;$�ȸm	��� ��F�������ܪL��^�eaN��BOQ|a �'�G\Q\AT9������Te�)8o��LNZRxσ�>�9�#(/h�!�/e!tg�n������0�,gvÙ��d����Ħ�i�C��&��S��M�܍��9���lc%!����P�)_9�G��֭ᢼ�f��L�Qy��VB�r��Ã!���g� ��UVE�������T_gs�J,x�%v./�ٟ��1�c�c]�'�:?�ݲ��K��ls�[J!�0��_�j�����v0�52�q�s��i�*��r���]�J*w���B��ُ��b�&س?��ם<���@p�L�.�fZrO�6�ͥ���*r)~Q�º?1^��7B�+M���KM���&`!�Z����=�ZjXAO���Q�Hj��~~ �-���"�*�	ķ�~�������qt��m�L���`�̟M�>A��Z�L��Gv����l#`кWS��u6*���T��Ha'�����	����c?FǤ7ބ��Z����8۩6�)��N�ӝ(�0�r��L�	4J�5R*���Ƃy��S/�X���Z�R�K�F��j7Om��-�"K@��C��űX3kS=��OY��1 ����2&GC�
R�:���~�́��B		�0B7S���
�Q��l��Vv���Nx�>�m(�Ǽ*��E%L������ՅX�6h�YŹ�:O��;¤����
�"��_��o�bju\y����Ξ�Y#����7G���K�N�跃C���8�Oc�%M��'@�E��(�'3C5g1O�8ވ&�~�LzR�!Գ>��Cx��a��]SY⛼�3���8fM�1�l֐9
��<u%Y˶I(��y(v�u�h�T!���(�%ͯ�?�xX`����r4��ZF*jMqo�G�\vٹ9�}&PSQ�:� ��J#pz��n��`�*�kd��!�V3WR�R�,gۉ�����%k�f5].Q�|�,�
��u+�����hƃ�=����.J�Z��;%+S�>������t�#L�"�8%�0Aq��C�B��D� �'T��\W[O�j�3�\��x��b�Y57��y�/[n��]gå���4-�JHB�y������x:�.�:el��d�����ݶ>��C:���^�gj���dT(5���5O���$o��TQo�?s#}����<"e�!\�	O�M�����DÜQ~Jh��r6�1ۤcK��e#N�,����Y��td�J���K���bqo�4[6�#��|�Kq8|�zV��a7jM4�yK��a��g�m�R�:NY{�e�k4b�܏1؃��#��!��W��@��o��5\:M+��U?��/"�ι�i�F�̇D��ȉ���wf�c�In/�:.�ư�;��їIU��6ge�-Ѝ��C�{�FoJ���8�X8���Jo6K]0�`ع3@}_ȏ��
3LW���te/�9Z�P$��힨s��`پ�4��7,��v-�,�[�K� [᤺���eUV�T��(@�,����<�Sۢv�أrg�m����� ���TF�����.\��?!僁Pj�Ie^|X�ܗ�&yꩯ�{m/O$z~��;���5A�a���Kd>�v��\���x��2���� ��>`���V�R�sLT����q�H���H�{
�s�+���mѿ�.���%��%[z��4�{rbg���B�2�ܰ��r��]� Zd������3�q���ٯ�:b�t��(
 Z��j<;u�� ����!m�L{���$3�bsD{�N(A|ϱ�CS�=}��M'<*h���!�zxZ�����A�G��c�W�`�+��y�� ����|��A��;�̵Z��)	��[o�S���E?�|�*�`#�~�݂��t��C�`��@��L��ɞN���b�!*Js�둜��^*́���9H%�Z��*���1���ϙ��}�)O\�gy\����}^�|+� )T9a��iUkC���}���c��^�y�u/qk�S�k)�����|7����ڟ�ت?Y�'Lu*��_jZ��6�ȨuR5]�W3�9���)<�h�D2��b�v"� (H�Tx�tx���?�*��7@�B�d��RX�{��em��PR�Z����P��*�x���$�*����ҹ�aξ� �7��N����䍵��i.CpF)=��$�>L$�w��ʐ������I˴�ex��m-�W��XL��/���\����E�s��z�'��N��0)Њ��ps���Z�w�=c<�:����V��X������kU\���4k�	�Dڋ��HvTx�术1�7�&QI��nA{����'�
���O���\�2�4��1���g|X�񧢰�(Dƪ��h��v����/��l�)��/b��Y��?��b�1��|&"k����C^]Vj�A�_%�]����F4���&�h������U[���l�tg���Q�<_t��!K�h \���&G��U\�@Q]p�6�%��L=l.@%�"j�
���Ʈ��z���D/*r�u�Żڄ/uʯ��F�xoҵ�@��|�̷Z�K��O������B�����[�h��}���֕�u��_����mO>�u�\ �	�&�_s�7D`{��JH�U��C�{��A��Kk1�_���i$gk��``�j�����Ԛ�9�J���-��&=�?��{v��r�mԔ��,�Tou!��W�QeN�[�N���8���	����\?���C�#���5����g�z�s"ɎM����vq���{�B��6�7/"rqq`�Y�������v���dĘߖS Q©s3�����6�~9��19�)�L�R�M�����}$2B����No�Ć�?��n�!p�.��9�������eUn܉��������d��Ң675 7p���(�i�pz"�����~��n}Hf�ɍ9�e�!Zw�^i�)�{�]��g ��a��۔�9�� �iA���P�����86�zMxN�����9>�9��M{A�SP�b�V�=\�]��M��;¶��Ұ�>P�hm���id���so�����k�,�S��рP��
C[�Q�A�q������Y���G�0��Vx_���o��[zm���7�(~P�Ru�[%T�5���.��{1�p�6���������t�5��u7��e��L#eπ��,X-��G��78�����pI�Z�=pz	���n��������'P��L8]Q+���{:�)m�Z�s�Aw,A�Վ�Qf� ��x lPս���K'�������kY�R<	S�����b��������b�����QI��ǉ �+_[|Y���M�ALd��8b��1�j���KD���EH),��g��v�vHzo�$�D��u|����{��s��� ;OZm��k)�J� {��
���p�;;�pl	qG$�a�e�����i�8�o��O)A�'Ζ)	v6`�P��q����c���ܵqSW�����K3�/�E��d��P�9�f7���5�9bD&!H��VrTA'�Mn���L�g���a��O5&�*Z�h������<����� ��~@���0�fCփ����V�Q]@	��6Nڷ	���9̺��hȩ�m�r9Y�.$��K�Ϙ�\M�>]7)�u<�!{5��Zwc�|E��LJS����^��GX���TP�H��B�iq����
�j�x���^+#t>��G��M����;!������m9�'� [n'�g�:S�g�MI~s.S�8Œ���_���kLB>_z'G���Ԥ��%l�~
55�Xf�D����:�`��5�����Á��wgV[��MS������Y�\�H ����\F�J7���d��Rj�h�k�ON� ��yˁ� ��G9�QV^�9�Ig{��O��B��O�A�Y���{o�v*�1��}q��5m��T#��v3�(=�VZ���0�G�$Ӣm:dg#�+ŝ�P�O���yFa���WC7�O[�7ﲾ��7� V.Z}�J8�0+j����H��ZZ�6Q4��.�ꬁ�'ˉ���֞��n���{BP�ҡ��]�!�A��_�� ��ͽ��p�`�Y�bԹ�AJJ��ؑj�òD�  Thu�dC��'o����f'��mH�t1�r�7�b/�zL�c���D��U����Tx��R�EU�N��ڔ�~e��P �����Pϱ�eU�;��$�����j����"Ȭ���E�C�L|�� 0)%����jCx�)\,ϴ�A�=5�'��'c�:)pS����J�&'9���0$O�{r��@�D�z>�yr7C���+FQjucq=�p���$��E�
�HA�*#�?��;z[�E�0����.��𤣵�g�7����ZI��$������p�y�����̥����X�xJl| f�����s�B��L���,!1���}������F+kثa�Q������������㿡�`ܨʍ��]WY��%�
� �e�f���[�L���^������}G�?��=�SX��^NB��P��,M��ZuTJ�5��|�L��lm�>9O:)X�M�����d����L7���^Ho,�-���f튎u�BgN��E��������
P���M~�2摸'�
�Acc��2� 9N����1!�� ��$9Ux�=�'�3�U�ӌ��S�aW.�,&�LY�P3�]H�A���.߱�ۢ��l�cW��z�tɍ��}\��/�M�d�P���yr��z�����{��cv!�qY�����?�"���?=�y$�H��j����̑Qa{t�u7�т�BZ�P�:�@xҲB����(��X�4�䎁����z?���S)S%��E���  �����@��E��Npw-;���:��:T�g>C�T��L˵�P:���p�M���#�]�F��)�sq�tE�ĺ�(��KXo�`
�[�a�:H��+��@P_b�" ���R�r�,�1�]s�4%�U����䈕k�Ed6d
�������#a~����çpl��Eڮ�\�vΌ#W�3_���C=F��G�@�h��z�>q��z��[�MeqP���J�|���C��.� �%n_�nA]�M�|S�~[C*�Zu\qS�:�<�����=J�#^�s�5G��z�O_g�.��flw�$�|k�<���q��	U��'[#����+m}.=��1��XI�p�����pC�S�)��ׁ��,�����]��Ӻa�r�,g���v�	������g���|j'p�)i�C:�hx����.(��`]��O����x�6��Tw��eWJ��r��`0e��9��c+�V�Փv\7q4�4�R��d���t�<�Z��˘���=��&,v=u���?��:�,�{x8���H��C��g@oJ����	4N������a�$�(*1V7wV8��X�.c�����R�-�&ܵ�'��". �[�#�4��χ�vH%���5������q`�<�S�bv�Sow61�]�j$p����3��e���7Qm�U��r���j-�o������"k�K9[�3fU���G��FP�"JW���I}m_�zjG����)'�:�im����h�6I7㔪z�Lx��F�J|�O�>�5��n/���J�c�ʐˌ|�.�Su]��$����-	rL���3����?Y��
e����7��κ���+�1��2�G���D�!YP/�(Y�ţa��BW(s��q���66U��v����%�aB4v�����+��$�9n��;kA̍Ij�������O��m�&�j+kc���c�nD���P|F�#x��&�@l��p��	���!�qi�}���5?�P�  N�����Cрb1[%��\�f��A*_�[���^]��=+$�3]��m���"벃"�s=ZU�<yd�i���4�5�%9>��n�Ѡ��Ҿg�Yfx��]��hX	в��/yN��:C�©�����o<s�O)�z<.H)�ѱT�R/��'�}���/�5��3�I��A��>to��H�J���|� 
�_>��G�q�����<��W��,X����.�d�ݠG|�z�����:L��dF�f�n�~��?H��#C�.Pe{�==���~��Q(�R�p���sU��{�#sK��@7�0A�}��O'����"����a�䭮���9��2�-���	�}:��g9����Gْ��M�J��v+����`�n�YE��H`+w�Qq_��`>�M�o4뙓���Fv'�:�4���nh㶭�`~Ş	�:hJ��?#҄���AL��D���Sv-�;��y^�������#�Jל�|����a�	�w���+�U�|��L�	qk�6tp�Կx����q]���f��j�miA(�&�s���P����{<�ć:|9E���j �KLo����)6ɏ�M�f����N���}�C�i�)	���b쓯9���z��b.�2�|C�g6��x�q�6���/��#>Ǭ���}�/=-�{�
�v����I�F/+$BQ���M�0�ZcB�g�.�kM!ḣ0�)Q� ��k�rg4���0���
��J򵹧DR�f�8�#Xz��-�?a�x,�~+<pY������>��	���莰!�iN9������ K�ۤ�nb��`JǷ�H/����k�V�h�lm�tf-�1�f�O4�%�B�1�z��8��5�*��3��m�Ngc�eɜQ��0�K񁖞8	�[N(�e���%�
?�����/+*��H�)=\�wz	����Jq��!*ndH퍟V���Hs��9$$JN�R��kw��}?��e&�W7�v����l�Y��=��~�9˯bz�2�7q�)���u ��!������k�&��c�UU��;��_l+�*.�?w����h�a���-��RSR{u�;����zH�L�!3�0	n�|���|d�r��n޴�.W��6� �:S���Z���k2�����}�<ٔ��-2yd��Ѧ>�����\�|�
�W��?R_�L����;	�Q��^�K��Fco�G"�f;9�1h.%�2�JGyF�Egr���^��Q~������j�v�R��zՈ�0č��<�����k�8��ǐ�I�O��A�>���O���&�Zy��E�m-�M���.8���P��(R�1���xZr����e@�2�h��x`V��?�R1�,��S��A�� ��~~��>{�A�ϝ��L�p�	��wʵIb*���$�����Xh7���8̝�μz�U��n��/����%�4�1�CQ��ڗż��/���(���M�?}Tln��:��&X��1�v�玸����vOq�=��IM�h6�ݥ �BM�����=N\2��]�~n�n���TO`�ܕ�%�� 5�d!���H�R����s��Jm���5���S�`��/��l]Í�������A�?�B1�#4��b���c�y��);��iT�h�۝NU{���*�>&�>�Tc���	0�]Yi��D#ja,&Z�f������R�]x��BIwf�v����`�up>���07Za� �ϛ�����ˀesE.Vg	�ʋ��z�a)���r���~*��c�2ؑOP{�<kJ0R�?î��Of}.�>�3��!�����	]�Kl�l=\xCy�1����͉&EG�$�S*��X�b�n�h�"���1�|����M(�w "[�kD���^��5���3U�3�!m5��fİ���/���2�;�ܣ����u��qԏ(�I}TC� ��t�������}.�!�W�ɣm��?M����OI�`�����ׂaV�>�Ǔ�c�P��h�{���5RFi�ÚU�NhAċ���^��#w�+��d�&���.�<N8x������A��#���̧izR��.��5n�]�� �	`��|[�vg���뛨rrگ�rZ��=�'���D��ϼ��!�P���X��BLU̵C�_k�6���,of1�G�� �"6�4}I{�r���d�y(~ �ނ����b�9@H�OQ���@G� ���q^9�3ǖ�/)\��î�a��~�դܑ.[9� ���#ܡ�Wq�	;��`�Ǭ2�>�2�H4�l��o�����Ș�uX
x����bŲ�c@�����_���!�4�dW���p��U�@�t`�;ZY�����N���N9�{
��VF�|��&H )�%�9C���wi-^�j��e����� ���,\�� �%�2���;$���W$-/s�a��N��=�S��/�D�y�v�5��I���=��&h3�_���7B^'{ǩ���q�qT9Tz�շ�!��o�ȼo:��Ϯ�vV���0��s�{����QS�e#�18��m����C��I��6���ၺ�j�M����lS[�����Ud���0i�3ݔ/w!Y���Y+#��jOʋ͠�.@_E��ŋ+�A��]D.�S�-ˣy6�ܿ�y7d;����`f���≢�N{͉�O)�����o9u��������]ټ��J���	Z�Ѓ*��H�dK���v�ϒ�4"�SdI4l���[�[���$�]���w���n\ L$���;k�i3������㶌�('�7Y*�xbq~�����M�Ka2ܓA�O��X�,̖���<9�X9˲������:���c��z�L�-��ƛ]�������0I犷b��s�DEQ�t����ڤ'�$=\��
�9>LT.�Ӯݶ�u�����YG���*�$��#=3i*��Ұ���(�`��K����m�)��S����0��FM5!P!���y���a�NJ۬��C��|]�}��,�4�e���f;Gۅ�X����,E����fzx^��3��$��ڡ�P��oOnk��)#l	zj�BI���%Uأ�?�{����!��t6 @!A��'UXk��S�O����-A>�5��-�۟����
���6 b���r���E�[d|���t��g�L$���#�5��J��SB�]Qn͉T�K���ɾδ�d�]s@-:��L�4���V�����T�ζ��iPY��9����ET�묢�v��B��K7��6m���V�Jô��e�7H7�;�gpl0 ��k�f<��+vH���ӱ��b��������sH�����_�;ό)S�\j�"|7����#�&������Gphj�r�`�L{턬c�&�\3��f���=>K֪���������V�9k�?�s�x��n&���)���*)|�Ǘy���?r���p�[2��t���D{O���+�_��1ُ���;Q?�E��̩��ջ�+�ױV�4�� �n#Ϣ�h��)'����yG�Q�l�[gaD'q�"�m���K�����225^���F�|�s`2��^�X��K~��@鎕ƁxW�4��K�WWr3YX�1< ���Lz"�]G�i���[m\̒\��߸��e��7��G��Z�r�����8}�*��.��E��rv`�W;t3%�x/�o��@����A����I�!����?�4�N5��dԍ�Ll����ڱ�Hr#�Ȝ2��%�"�͔	���J@Ex�SŴP����ܠc��Lx9uE��>�Ŀ��S6���:h<��f��a��{��l���J�b��(}���{MB����M'���K~![.���HP  ���=i��i��Ĉ�nU�X��̤E{c[<<
�o������x��_�.�j�`�w[8�VW�]$j��!,D�?��m%�h��d=�sK^zG�<�U�p׿��`�@�f����Ty�6 ��9��AUd�6>s�s	�OʠeD����	��ln"k�*�3�,�����nhX�i`�@n��͵"�ƆX�& ���0�û�5w��rD���oa)K߼��`�Hp��8	Y����4:�!��������_�ϥ[����ӸE[�uL�L�ι	,[	[�ˮh�I��o-}7��'0�\��C!�g��Guu�0>�Ʉ�]I(��kn��0m0>�y�HS��Zb�J*1B�,��1{���yĵ��.����L����Y�FE�q�m�讄��3'w�V����sjM��<��4���X6�� *��s<��d+��Ve���݉��l���q:9_Vd?=b_�f�!�@��e0 �_�}4b���k!����,;��X����X���<�7��=`ܤ_P����!lQ��:w�L��%�d�:<~z?��O
V<g���1�5#1��(B[�k��x]=-y(W��a���G��(�؈ē/T"`#�f�\���#�@/�׉@�#�ޔ���B-��H��W4�M��5���_U��ʩ�s��$�w⪾����(����v��~���.�_�9��zZ^���O�8�vg�*Ȝu�+ \;��:6��m�"�|�]�X���ܲ�ԫ��#K�B�=�d,�h��C�;]H�a�hE"��T|��i:�]��u�N>\ \���pY44�����M:��Ð��K`�43"&����>+�Ƨ���X=�}��[	;�u�W�����ȧ5�p�l�ޗ���+�����]�7o�{_dI`��!xHil�	�
�ץ]�D5�LR�K��),5]
jS�K�A�(�٦1{�t5��w�b!d���~ըX¨<1�P��E�T�W�\z<p�Ԭ|!�z��77BEf��fݎ��1�5��N6��qƸ�n��qh�g�y\�BVZ�{CָM��:پR�B��|��P��V�:��7����?��0Kx���G�
�U��3���v�"sf(l_ti\$?��,u�9�" ��(�s`�'f��&�y�w�c3��O�pP�[��@X*N5�����A�w#�\�u��䟁 �|���~:F$��=Ϧ�U�C��Ӫ�@���ml�6��qpJz{��7����P�<2���T]<�@y���-�s!q�`y⊚�'��[��/*_?Eel)�6_��0U�f;G�J�s��e�#Bիc��99SD\�5�p6R��M-��@�,Y����1]����8
�>�<|U���Qd�P.Á���0e׮x�B�ر
�6���B�&�kǾ��>�!9���=�c�횯���އ�O��c�	=��F�~��i�U|7'�{���]l��@A�b�A>�p����}ہL�P�N�QǏ�o� �ص�!B�r��,a����Er�� ���λ�v�i{A�}�}h��xlM��b�����B�~]A�m��2�<��VJ%ocL��C}�����SƵ���{�}x���6;0+�q2��89yj���)<3X<`�>�Q\DiзA����������H/��u��Dp>?T�q1�H�+�(E��C<�d�E�ͰED��p ���O�Q0�Q�6jڎ-ӟdWBzT���dlY��n��@\�m����m܅�u��W��:#ٟ�.��Ĺ�>��gJZM���^ӻ���vP����P��"b=IZC霄�?�)ۻcp�)����b�+�n�Y�[K8���K���q��z���,)������9`�uk��*XHFs
� ��g��X4}~A��;�J:s�:ǣ� _&�9#��=�!ψ#�g�J��b����4���	���#Ƒڄ����֟������*�p+��Eإ�\��d�:Eh�װHV7x���s�����I�ZZv�#2R�n�<���M,�ª��>.:=�g�~G�e��Q�5��}��K���tJ�*�_kR0� �)����Đ9:+�h+a1�M��ބ��H�ѿ1��Q�(;87��w��O�]�J�p1��	$�jp�
�E�[r��Y�6ꍍ��!À���Fy��UI�8*}��W��P!����F�橃=B� �}�%��b��{�3`V�py�܇���+Xj@��LO��O��C���s�d�U��g@h���[<(�����7�طxS�MZ���FbP�w�I-��筵X-h�b��Z���Z�k��~��ݭ\ O����m��.�<�,#�!�Ҏv�#բҫ�� H7�$�fP�pg9��P��2ڮ��Qd)v�%��x���b��ͦ��d�U�uSd�P�<b;���C{.����A�qh��A�'8����P��Ev�x�tqe���m�<��4����8�lQ��/�(���R|�7� �	N���̱1�C������/_=�lku�L�<k97F��fTm�����a�;F�P8������_N<3��3 	z*����0j��Z�5��i��Rh1�n���ؘ<9$�mDj
�d|N�{UU��F�[�
�؛K��iF���ѼYݺ�&b d�1�y��P�;��6��=mQfp�qWªBĚ��������@���h�ς7�q��3܃��щjm"�[�C����p�6�U�{��㽫(��}}����*f���Zi���1�D䮠C_��Ėd�JT��R���*y���'��������7Y��ڨD��V�a�g�`^�_WVn=g�!9Z�|�?Q�)���[��e%�b�1VT�������l��z�6��+�&eY�H�f��lB�C]��dA�Y3w�5x�����>}���G$�M�m�=�l�&�u�Efs�^��O��`&�&X�u5�)��� (�JPY�xL�j^�h��Ĭ��-���ܜ^yʠ����%��k�?�P+!� t�Y�TR�	2�G��i71�w3̦DE�J�>�ɜ�D[$�K�u�:˻{�}7/���h�Ͽ�u����o�U���$����@?���*)��)��R�]��d���7h[�%��vS~{��4h�������������|0R΂P�8���֧.�j���ҳ@���v�`3��y������;s�γ�SeB�H�J�}֞���I��ZO�f���U/QB���N�Re*fr�c��5�X����p9�3E�!�R'��v��+�j	 %y�	)��SG$�����1K��ѡ�.k��I̧���R��OE
�������aNR���ao7�!�9���v�j�K�i*l�E��*H�\��|��<�����HC��6A�|�V��b�u��!c�F�e�0�電�Ձ_���[p�Z �^9�y����q��:"��Ob�N�չ+۶u_���)C=��1�zqv&f�LH"a��p�a/cLHŖ=Q��]w���������F�i�X]/��6��u��ɂ�4y�J��z���d�/�I�.�S"i���BE���h��G��1����2���Y�֩��c�vڲ�o�L��/����'��
2>J��`Ɂ���ݏ��"�~%ՖO�����E�}8���He^�����&��z���qLj��4�Ą&r��D;tU�G"^nr��v�r��t�կ��*�Eb�i,��ZZ���.��đ����h� �`��P��i�u蘼��t{ �GΦ�4 ��P*|fgߋV=D~�T��]N�����JD��]f��@����U ��d�8L����f�чq������?����3.:�qٓ�|�p]S�%�����S��n�Zp�.X@�q���.oS�����BIIX���>,�|<�F9��E��'X� ��U�K=~����&�D^���~p�O���I��׊��]�'�]=HW�$S$������4m�PT�}��ˤo4s%���z�VDH'�'�3�0��a��l�Xi�f$�P���*�~|�$����UP̰:�`-��r�w� o���"��d�2�(h���}��oFi�uiV+�A&� �H|�A-�mӭ�&�.��e[�s��O_vW5^9��.���l�h�s�*p�[BR�FF��Y���$�w���B��]>4f���,w��:Y�&zqI8Z�G1.(}��~�l�(<(Q���c�]�da#�W�(#%�C9��$Q��r;�������83m,[C8orp.��tn�h*?�>y���%�2��Ɉ`�Qj�?�[*��ƼĢ�&nT�Z���z㊪�KZ3l���R�����M#M'_�/��`�� �\bZ���%�z��ǲfu�MVS`�ѓ7��"=����(+BY���Lb29��(���TI�m��!����h��NjH�
�=^%���"
�J���A�w���p��J^��@��P�-j�wF�mx�s�K�;]fЏD~�}�	��/��dM
�*��D���L[��>��n���*���"7-��+��qR�_��P��g�F��G������>$�"�[��ʠ��bD�a&��]�ܔ��p��7��)�F�O�N�%�ol��h���O����8�ZX�q�EkQ0�$`���D�������w��NA6ʍhy8�Zb��H�^/��m<�c���,�mٗ>
r��p����]>noG���N�ϭ:�[�+N#���pj>��L[,?[Q�����'9��p�)�h��������m�-���vÿT�āF���$���Š��>���C�&?^�����+S��¦��- M�K�U���}�����n���Ε	M=�
�N� !��M"1�����M=�1��sFn� /J(�';�v�i�6�5�%^ᴰ<�����,/��yɰ��p*��X�(3����+�6�}TB7��/Q���"���Jx�?��qC|3K��Y�u�IO_Ɗ���rOǪ��FaJ2���OW�쒄��!�<4f�D,�q4�ؙr�Zmc�c��e���a�(^�6q��fLX�X�z�Ř�B}x�p��e�������k>=��+Q�^?���90�s:�?�*oG�͂i]n1ܟC�����	+a�DDᢖ��#d��IڥK��tNR��004�w]h!30�l��i�߬���0�ɋ��a`C������Mi��B�;��
�9�
�����K  �*�]��LZM�QIZ���97;_��,l5��A��U*qJt��!��籇�ċԈOږ^���r��C9�;��I�W��� ���F����~�!a��d����r!�;s��C�a��=_}�5=�����Ο��wi��(��b���C�;A�6�#^5�W㷐CzC�:KXt!a1yV�d��S��	6��j�$X�j��c��ŧE�m��#�,Nz*�A'�R�y5X����[�:����+�2��	#Y<7��@��^%FOS�44,pt�������h㣐!���n�B���VBҞ;1n~:e|`r5i�yu-SME�t��b�4�H7>�X)��ʜ��XJ%|W2ظ@�/7V��5E��OZ1�=��Ĥ���������xW��³=�0S@0�%�'�_#Ձ���v���K��y��M���sy�_]�|[�����(?��=��L�[�Q�Sϋ��P���][_h
�TM�\*s1�j�A�_|��C��ڳ;���0m7p�T�\�wAo��R��X[6�ՙT�d��Î 6a�w+����z��q"��є¯��^UԞ�|�u[ߠ��+P��c�2-|���/��f{���V� -�L��_�b}ɫ�A�B�Jrī����7T�
)ɏX��K��3�,z��1դ����啞3�o��##�����
:�q�\����j)�N}S�.�oee̴�Ǖ�FW;V�B�9��ܘ����K^x��>���������a���+pUC����Q�k��r��n�����;]	��h����3[�uQ� �~A�a��WARj�x�����ׇ_�]Ex(����oϩ�%Ӗ�toD[ʻf��=�&w����mB��Z�Oٵ^K�>��<ۍ��X$x`�A��D��S�Þvv���ޑC�33�$���)�%)�p��Lpb�8����G��LP�}*g$�	9�(w||>��^���[	�?��t��<��Z��M���^HYhdbd�*L�è���M��Ų�~��yrH)@�Yd�ry��g��T��<?��rG�s&��z�r�vi��DE]��pG��f���V�!���$82��?�v
c�1���<��o�O��m0��lZ1X��f�1��I1?@O;އ��f�<1��'q��{��?�P�r�\���qN�0�@-G9r�
��j҈�t> �5��ʯ���'p�m����e>MH��g��'#B��6NP��c=���#L�k�d�j�B��B;�H��,���|�4�����j�'ZZXx�����J�{�6s㚢[��wS�KLR��dn���+��B��|*���g:���xvS�ch}$b~L�B��)O�;c�_�b���L ���8�O��8�q�_��A�_�Hĺ?h�L�����	����f��$���{�:B�:��i��"C�j~T�{?�6yVs��6e��
#$�E�2R5n�f➠��rmæ�:W�RY;���W�10�8�/J�n�V%��O{i���pf@o���t����	�-��T3*�A�����P
��/�e�����۱���������az�UX�\��{F��9d?��P��q�����`ϣ���}��ӱH� ^V��YiW���g!���cI��2p�cCN�� N�=t��Oݺ^!���5�Py����e޼y��`����`��iԟ�1�@N��۩_�4�i.��EJ�&X1��F�� A�͹/)$u<��798&��%J������"}:����*Z�"�Q��Ź�$���?l�W��2�'ؙ$��'�-|�ѯ!�a�Fw2�xvﻅn�Wi�FD)�3c+x@-�<�������u�	K��ɽ��JM�3��l�P/f�CwQ3�:F�.�Y����]�>it1f6V�r O2�:�e��ˣ�?�\.Ͽ���8��� �d�u��/c��<iNZ��f����s�rt�_�o����n��{i�])6�-B����čR��ɦ��-C2�#��Py�I�/�ߙQҏ$�q"T� �`�@0����6*cv��VK��6�����k.'�e�<�XX9�-�Q��}�#9G$�M�}�� U\]���_�S���\)��C��L+���W���p�/�[1��r�q�4P)������5;2�X�	�P�P/ӈ5q&;�9�.b@zG変&6Ѡ��3o��J\�͡{YS\j�I��f�k�)`b��v�*GX�ͻY�F�f9jH��oX���;�D>"b�I�h\y9��`F��6͗}$�c�F���Y�U����9�F���p^܇��[VԾʥ������f��ų�e�ߔ��C.qX��83��>�,":)�e/ *�5��},;A�4y�E��s�B���a����б��x���h�i�	e+�]j�h6��&IY��;7�'z�^_�W�!ޓϟ@�F�b[Ǩ�K>�׶���� sk�Im�/iA�D�!�0uרgɋ���sŨ�uwh
�3�x}~ >�w�����8uH��E��ђ�h����h��х�{vz�&xUчUw��31���g|m�<���
R��W�h�t�ܖ�>y�vI��J�3����	���'�7�'�������Qڵ�b�AXW��כ��X�I���#"w�*��T(��V��.ӧ�@#�H�$����s/\7�z48�G�9�v��uA�h�Kp�=��4��fF�N���.<^~`.�����8͡�����)~�������ݓ������>F�LdV'�̆��(��Ԛ��z�w�LCc���.�90�6�	&� ��ȗij�W��*[�5��4��nn�q�hx��j/r*�(�r����m����\��'��X���X�!���_ƫ�Hҍ�1�h`�ھj%y,S"��U���ǂD�0d��̷�Cz���œ�W���BŽN�kҜ�}?8k_æ���B�R�ֈ|�v�/T����u�5��T��y�SM�-��[�HZ�%�ñQLm0Z%�i���cI0�� D����-�z-5I@u*k}�O�E'�t�1jZ=����`́[ٷ^�S�ys��ѝ0H̬�� 3뀼J���7\my3��,'DX�/�����I�*�ԝJ��ڭ'x������K����u�2~seˋ��@�,C:hZ��O��p#$b�� �9�v�9$
����7���dѶP�@k�[r�y���?��p��5b4!8C����>}'d��c���X����F�����}O�<��!�<�:��od�M X�.k�
-�zzV������JA��DL������RQ5i�;�@*�3�*�Y�9ڑ
�Lu�1�S�S	
�I����!�� �n,�/kp�?y�o-U�;5��u����e�x_�e���\�e�y&&~���nn�	�d����$S?�H���"S��rPR��9�BR����;�e"KYhٷ�O��Ӏ�O����ap喩B�͖BSB���Wx~�b����D�#A���|����d�\�h8�:�ݧ��	N�-����]9�8<�bK6��+��@!��O�੾	w� �@�s�s�&��׺o���r_�8�m�}9�������+Nj<}3�&�*��1#mϞ��oXoPj�֬�{�������ۨ=2��7`�5�j��tO^�\:A�A���͕���Y�P�����T�{<�[�@A�\��$J�W�^�0�a-���qq�AX�x%M�>��hKU9v�K�|H�)���y�Ӓ�}	䝨=s���QU� wP"�a�Z�8��^���Ġĥ�C;�;�����(���0ɫ��{�y�پ]F�����?����v7I����'�&Rφ+����W�;sM����\��m;p1M&�I�o%���o1Y�_�7yHx�';�U�8&.b@=-�?qf2oψ3��P[Iy�u��^p)��t�^���d�s�r:�N��<ڕ�8$>�H�b�iL�P8�J)���n��bMA�UD�{�pSs�BЮ�_�օ�2j�H������2]�'��&�7�m�b�	U�����H�u���&�?a� ��U�X���ݙ)��r"�	����ME֏왚��4P9:��s����ab?�{��$�n��T�Z1+���,�� s��(� �\7��n��|#�����n��aJ�]/+Q�L��;%6	K�B���{&x�^�x����{NV�:��a�z���Q�z�(�e���hݤN�IWf�Ao�.*���SM+�����Ϣ��<��b��v����G��5T;42N��q�02�]��m*[I4Lkι�L��]�P��Cg����9��k��t�[Jz&��\[�d�]�o����d/n�E�(��&�/mЪG�oWM�F�P�c��o��mA�մ�AeT��]W5�	f젚�m�����)H@�����#Xw�T�r�mh�kJ?�;��φ'��߃��D`��%�ͤ�����^��M��!�UF����b$�&�_��"3T�@"-ޜ�V���u�Ic�]�}���v9���ʍ'p&U�8����g_��ŗ�%5Z�$cUb-�(ь��r#7�a���KL~�w��'ݱ��c��A���#lkO$��cU4<o�}n	e�`QF���;o>g-�]�H�
nN��b�P`馤���*M?����{�ZU�K���ʤ���D�脰����ϸ�T��F ]�z��K��@�pgv�!a��X��WQ-�uF�2xH�6#l1o`c�q���1�Y\)����	h�Dm�AHq�¬���n�t��*`G{���%1�:���V��6D)lmX)c�C]ω'0yOe]Ï��^
�x��h�
�)�`:��?�&�ο���$���[Q}�W�h����54 (��2OW$m��{[Z�+���E|y\��$���*�]�
���~V!v<��x��\6UؒK���ZX�O�l�3re_H+[�� >�`�����=�LR�z$��}��I`#$1�,�۝��)�%�p���񲥨րo�d�z��A]�f�R�!�A���4H���gO�g�&z�S��B���ѭK���KU79{\��h�y&����&�h���#JӀC��.���`Nx�$K��&s�h/\/b�˘��|�|0�[��M�&�xSG��%(J؊�l��2R���i|fV*$V4ڔDz��\]mDiy�mۙ��	.'�2�3��c�L!�U b�.)��%��-vU��L<���;V�{U/b�!�_i��,o�v¤�b�
|E���3�{R��Lvp/���Q=��*�<v6#�cb�\�>��oSP9��{�,t�n83������qzE��[�v��i���*kg��%nG��r���+|�Jp�t� ���7��)
��zMXZqv�Z!X��ߋ9�e�P�8��	&�t%.H��@�O���U�����h��O���7,Ԍ��;��x�p��E�HV�)��������@���iTOyAV�h#�A�_�ʶ������m=,�$e/�?u3��2�����a�U��Jn*XW̖��g�E<������FF�F࿡�?��H[�<%½փ~;�V�%�G�8��|������tHa�[E�<�PY�W��ʬ��TwjJ�f7,LO��u�����(#��!����J������sv�>:�E\�ۋ�^W�3��3��}�y��c7��B"_�O���1�нď˯nDSSz�2�(}�E6���Ѷ<���s�N�2OB0��x^CFOt�o��}A��z|7Á��9ץ�#^��`2[�~�����=.���v���	���fፚE��(kU�5���m�Q|U��k��	�9k.<�T�:�,�sω��-LQ,�6ά�s�Xy ��.c]�OKG��DAE�����Z2�q�;��)AJU�S����;�lDv�`��J�2�a�~��f ����}Y��uMB'�p��&)e�2m�p�z][�Fr��,R={]:�]�e����YQ����+^ ��2PN�`qn&���K����)�PjeR��ӳ�麔��o��b�����4��Bk|�z��t�Z9�n��ϔE����ʜAB:d��\��E �%0�BKè��=���e�4���K�臑KTL�f�i��^>��hT�s�f������d�M}����,7C�I�AY#�>��^�׭�#�����'��fʦ�G�F��W�V2��"��M���8�˼!F�S�fpO�R#�ƻq#n�a}c��.g*�NѸ����%� �B����;�����?=��ظ|d2���+3T,K�~
'�S,ǎ�
��Cɱ�x�� ���[T�+湘��˲uش(x�qh9Z8��C�F^�G�E�'��a��[��u�VSJ
��X��+Ǧ�jM5i�7K����KN��X(��FЇ������<(35��6
M���b&�C���%6�/��g��;'f��	)� ������U텵YGE��hV!�f�fgGr3vgj�����jD^~�����e��9�|�>AĎ��.k�L@����^�a�p��Z4�3�5�TV�X|I��G�g`!]���J=�	�����8�@���h�Cص��`��7�lU5����$�u3�>� �O�[�����:H���X�tk#ّi?EQ���'&�8�X*&�x&�[��>���vձ�?�w���k �P�Di�}�d�<��+K���즫��l�I��I�J"�_Ph~��I�]�2���8�Q%}|���И�6�G`jm��΢�����0�[��#���b �m�Լ�&qɰ��#����@0Gc�� ��z��i�H��h�_&4�����R"מ��cK-厤L�:f�
q7�re��y����^zF-�)= %�Xx`����vZ$Ci�=p+��,��P�rP��J�L�/��g�����P�B�mz:;�����LU?ow��Q%� 7�ˑ��ޖ�k���9�F��P�1�կ���F���`ݴQ�r7�B�������i�(Q�-T�Q�=H���'�4��I:c�m��az	�x"������lA�`+�����C�V���A49��ց(��3LH*�a��,��$Ѭ������4�VD�Q:�ٴ�&�8��A��To��0��,:a���E�<3�w����;�/��teD�`�6�Og�|�r���f\u�ʺ�֠���o��#��K�mT�ژ�F�qج�sKƷᨽ:z��X��Iɨ��?��V������Ы��cYqʃ��ON�'Sӕ�=�1Y��oE������S{ ��T�i□~B6�<h�\XY;W��5������-�X����{���h捂q���]U֠�����c&�vZ��b�S�ҽ��)$�U��9|���^��:m8`&L�.����;t_.���@mn�XA�{��g~�w���Up���
�
�Sl�f)�b�)dK[깷7S4�zxr��eu��8�7�_"��ŕ�^�r�-*DWe�8+&j&�f��J�X$}�4�D��yY[=X�5EAL�+QBůE����� ����.pF��8w=+�,���졛
��w�t�C�9=�fW�|5
!�hk��nD'�O�����Y��kѼ�*ƀdT5 ��lN\1i畜��뿢�
!��*��)"I�	�$��k@�u[�5^���{��ɪ6�s�U�^l�w+ѡ��&��g^�� J�~@a�~,��#7!���W�|�.h�-s�˙�>bS.��)�L�N��w$����V54XI�c�I���!�8K�rxa|��=9#vL��-�J4��׍��`Z�~y}��XMA��u5V��\��iGs"2���%-���|Tl].Sz�a��[Ã����������4X�˷ :������,�hYZn(�����.I��y�`A��]�@��t���ŭކ����Ji�����Y��ǧ��k�u�>��_'���S���L��u;$�:���oB�~�Q �	}ֲ��k�t1�j�6>V��1^�̲*�YZ��,�Z���n%ë���)���{��UCM�����M�^z���T��-H�,��Yi5��S�e^�9��տZp�d���k�sm ;��Ybø���X}�X�!�������e��=��P{)O�j�,+^���BG��L�\wُ�԰��ĭM�x�ã����Qȶ+�r�A��gg�)�3��X��R^DCf�f���MwcA�0�Υ��a�o]m����ƊmXI�>^2�_�,;�&�IW��qZ�Ee8U���r�tJE@�Br�f��`Zf}?@����� �|ƺ�	�֑&�pt������/�Ë�s2�����P�J[�����p�D�*~�f~��$o�r�6v�Z�?Z����6��>�N?��
���"�yc�ϗM=�`" k]U�V�(� �/�#$�}ɻQ��p��Eg��� ��Kd�!�D�����__C!��1ђs���v`�Y�5>X9->]|e3d������y�ma���T�N��8F�ΰW
NL`h��^��M��Т}y��́ze�9�A�9 r�2 O��i,����'O�1�D ����g� p�\u���)ԛ&�аz*�s�[Ȅ׊��lZ��+����z�Uـ�Ɩ؊T�Uy���U�a�������~�P_�''<`��j��3Z��*g��Iy������ܻ��	��t�~�H>ǞV"�ΈX�e�S��Vz[:�kb���r�;�NNZ��(�2|GT"��{���@Xwr��[]j��J�E�N�q�@1a��iV���j��K��)�*=l����C _$?�mWD�zʘ �7/�����jN�p�M����ɤ����ќ�r�վ~D��M��QSeD~ ��bč�e�������+�v���� �'�+�d�]ێʅ�}DBz3IDyd�8t�:��$�r̸Ȣ�U����5��"�B�R��Kc���O�/J��<˄c�	�J�
A�O�N��(�(eP���^]�h��o>�g����([P�������[jyakW#�����P��%%�=Ą{�Y �H�� ��n�<��\�6����Q^r��и��͑ێaQ��V2��fUa�4���-:k��� ](�n�Qo�4(P��Q)�	F0�n3Ô[(	
�����*�},j�M���?���I���N���5�È�~a���
.�hr��`KۛbOs�[���C���Ǔ�e����!���VyiڋþG���q����{���2�R�>�ݢ	��Pl} ���h�e�&[<%��ugCz�zl#�oP�Xb�FG67'���J"�ox��=���DŴ1(P>p@4E#,�)��2%�N\m1�S�}���p��~ M�}8�8�����ӳ�!�9%�~l�P̦ߠ���
���!�ʊ�ØC�m{�"��p�Ȇ ��ދc�������iƔ~Ĵ��zY+h�ׯ�{�W��9x���"�'�:�E����s�	��>�����O'��D�wx��z��whN~{�}6H��/�w��y�_ ��hG,B�@�fDj�G���T�>�R(dVm}�<pZ��᱾��6��^ݠ4㝑�u��?���f����v� L#V�xR�m$Ջߍ�#R�{�15�"�Bȿb�u�� ݽ��#�`0�?t����ɿ�Zz��)Y���\|���
�Q>�i�4�ϮZt1j�� �ݚ���C�];�����)4g��qx>�1T��яR�vHrBZsx^�B,�R�xrF���������dh33s��G[\~�]6� ��)iM��(�������������RR
������&��|�c\�e�J51�����i�8�Ei,�@Xc�c`�"<�9���'�w��c��٭#r�_�؇��� ~!�����Ԏ(1�y�,*��䃁]k0&9�s��mR�����q˿��;���J�T�q�%S��6��;x�ʝ�\���:@f���/ݶzG�c*(?S9�Z���h$��y/m��@�%������)���Η��~�#�Hp�u�]�(�C�Xv��a������;���/uA�wt��r����P���I^�M}n2P�l�ݵ�`H�؂Q�0!�f5�	�l�KZI�b29��~�3t��R<��"��C$0Ze����rKI���3�K�*�$�)�
$1�}x���Nq���v?���	j�����I��v+��4ܢ�����%ry�#�|�ke��)D~�~[X�Gq�%ݧ�豔#W���*����<��ì[�`��М��Nyj#�	h�o�M��	��^^��7��O�=��Y����1]-�2H�	qO���E��V��J y��q�+?�C���O��j�_Ъ�5q��?km���B��C^X�b"Y_�v�"`����	�a #�Au=M�im2M��خ w�ُC��
2���l����
x�8O�	�?>ՐA.k�淊���A��x�L�_��(/\AJ�<� Z�O�'3�p|_���=�A��u}r	H9<��ډ3t�wp���� C��+�=������'
�u3��F��,Sb����7��-��W"z��Of���A7�`������\Mr ����v�K]�oͶ�G���F�ZaR畦po�����8��?����}~& ����4��],`�g7�e�8��,>���K ��աNM�MI��ZO��"��|1~��mxe�]7g9 ��1�=���c�t�����q�<��V��D�oDn�<��`&/�2[׍���e�zb�"�"T�XH�I1���m�6�E%XC���˘�-�EvO�x���2"X������G�,����q���@����8;����	T�mv��e;�is�r3����_���w��[V$r�G�W��X�f�%/ZSf����-VZp��k��EE�pg��@�"���h�R,�>����#�&���w����K�U��=�\i`\�\h�����G��~�^ y3S�S� �t�a�>�A���H��Ca�bu��2A��\�I���Ð�9���? `��6�zcS��:�dPw�N�w\���H4Y*��1ZBS�e5�
m	'3��@wrI�n�̞�e�Q)8N+� �]����wS�b�|9q�x
,~��@8|��y�R?0�Ru�~��%KcoR%$cޮ���(|�.B8\w�}'��X`�s2�;'@�	�=�F���L~S��p�� �39��=�,g��#��a�`��I��Q�z��X�� ���v����_�Ո�Z�Xn�q��g��h+����޳ʣ)C�/:&�b�u.d]�qQ$�JeZ0�i\�?�C�οx��{��k�6=��.Y:S�m�r�>���~eg _;�WG B�;Og>*m���j+ s!�A$,�J�ɜ�lK����⣦6k�����%�ܟ$&3t�ü�5�:%��U��c����Ɖ�ڴܹLe)�p?�����D:Ê�_��6�(>l%W�S�.hEfs��DG��B�s8����ݣo���;D�g]gQ��f�_��ބ��Y#s|mv��N�����k�m����J
��<�� �5�NT
 >�bڛ���
kl���m8��SD�"����O�F���2����./�]A�a�5�t�fI�)��'	)�T�\����%~^�)��(��*~�YxʇEQf薍_�i�K?�rCm�b3iamg�jDr��W-Ґw���xzc8ވ|� �;�)�R9v�R����?c������<)�:t.�H"�ww}�.��=� �dV�f�H߀��T��D�L��7���T�I�`���m�? �}i��5���F�m�J{���,RЮ��z=�ނ��4uG�4h������	�M4����{_����h�O�\��y叻o�� �T�%� �'���綰Ck��>3��6����op�X�UKW���n9��u���P�uV���/H*p��Y��Q�LU=х�)"Yal���?I����n����M�e�Rl	��|��; مY�o�*�(��V
��v�<�������7%��<7��%j��.�;�Ln�)�2dJD�m�JNr��q�N`I�-R�h��i� %�*a7a��b������-�OÍ���"m�J���������\���WR�q�EfQ
�l���']?�ߩ��g$)n�Ww�br_�b[ur���(.��R!���޾�8�����ћu]�l
�6��S�a��J5�~�D����H�y�/!�{T�$�^�d�g�qM-�)�qi��tkm~�2�;�ƹ8 �x���3=�,� ��,�/W��]koD,ݟ�6š��0���S�B��I)�%�"�ѹ�{ARXZD/c�
�ܰ�_)�#�U�j��]X��,��_ֱ�4��Ή�LX��hrQ�O"0� �n�N>��?W�[��뜣��*�0�^�]�$��a�@;nH
|I��%�%���Ƨ�����꽲}׸u\ad�EF�������t��5Ƣ�P���Z>�T�R7��k$�/B����l���7���	��:q�����dO��n�p�<u3,�O-|�����_�w�{!���mq��Xp�0�����/<���5
 �n����¸�����`����Z'@�S��B��F���oa�!���[/��K�D3�>/L��P,�,6rH?%���5o��n���"���Ce�Vi����+��]�n�.�E�;Q��Q.+m���v�� )�~��ogZ�\�_br�
�5eU3|1�4y���ܡ����X�z��g�]$91�`�бJ��iV��a�sp��_��e���.�����p�g߿͜�T�������m
����B��w�ۋ91j3��Y�}VC���fI�z���)FC�	&�K���������q�^ˮ�i�g#9_��x;�H�Ly�����M��_��tfz������ �O]?���LD�����=��Z9_s���5��|�VN-���JT/,o�D���έO�=A I<��OÿGwXy�3�>��@s�����N&��?й��gn>�v�i2u��T�9�0�-:kkK� �~s�gD� _s9�-w�y����؛ ���|�e^���Q��@�c��G�P��K)\�� �1!!��3�r�Bq0u
$�9I��ڄ6}{�H0`f_�M�e���G�R�˺S��ɕ˦/&���f��T�r�T�hQ]��P�����TjȆ��#nY�SsB�a�/bx-S�5ݼh+L�L�eփ,�~�^x����'����PGw���H�.턑��:��1�3�
Ǭ/�\W֪;K!��+������<׸����%q�3�Y�.���T��a�Ӱ.ԣG���ρ�"	�/�kp�	T �'.����ez|�X
9�M������ߡ�COA�XyY;or�#��&*z��Z�t��	kN$j�ڛ��q�SL�:=�"�rD���bP�(��Ol��c*y����9p�����V�'�z295t����=��ћ�b)���}���q��<�c�=QpH� ֈ�U��¹�gBagT�F��Z�zӘifg�D��Q�����಩L�f�8�V���ٖ	u�r4�V��z_��X���
yXʱ2�4�t�I�u��R�g�d��y
#����}�>���#�u����|*pS��i^kX`� �K�欬X�2���K�x�/UP�����Q�����,��`�Rnk����a�$�L�IGt`������3�e���XU���kf�Y�Z�D�M<V�7aO@�b6��e�i{Ǣ����I�N��/��?��P��k[m�N	Qt�]���Fk �Hߐ�,�$����W��y�m��� ��`Din��_{/��Ǥ�n�����XP�b�,E���hkO��X����3�P�݃����H�m�R0���7��_�]��ۡY�U��$�e�!&�D�kœ���p�M?�����8��KI��)2�r�q�����_�jPq�<�r�*&�\�V��X���Y�:K��is�p	{.e|~:����7��	u�G��t�мJ����ň�����"��X���>���rl��g�>V�{��ք��r��"u�h$�Y발�u�RP�Z�}��u��q��v�����[���\����
�+ٞ�z����:Q/�����*^70p���2NA���� ���k�]`�D)���#*yF�O���ð�l/�'� ?�aa��m�P�[�qS��I�9s��Y�5��V}�~L
�>'Q�<^��F��5��/L�+J@�8�w&�c˷�q�\� �,չ�|Jc�2nBյ��"�NĿ�u\}����#ȶv���z�x���ݘ�i��}�%oߣ���5ɥ����s����:zj�D&���`?B�4�:��L]��@��4�z��{�s�~gv�`�����&�?*��8�J���r��l  �=yq���/'�'�;��b@��V�����x��>gu �!���$�i�X"�/X�~�:d;ڷ�c}�����GǇj���O㡘����`�6v��4�G{�ǲ��8Q���(��M����zʾD�"��;6lA�a<��(�������S#��Þ�'��9�v=�c�3����cc�q%��ۄV=��qa���T�����%��V�%R�YG��W�n��������pu�+q�Iq�׫|B[`f�"�'��ˀ/������D+#�0�����j?:V^�"�[`o��~���p�b�(w��d��ȴK߃�aq'�4>M�O7��H^�΃��M���3�+��G��)&�/�Uj e=D4�$�w{g�k�>��!L�N��ΰ	��2N����Ag�iw9�Bu:�����LMw�&���aN�a�S�dAΔ�PZ��l��L���Q6*���yZ�l�����U��X=�iz�G$2w]7v	��n���ԉ�\��{S힛���t�^���l؇�8�L�	~*Di������O�䟉u��/ ��)J"4[��/`X����s>�G�fa��q��ܿ-3�h��!���h^��b,�`j��璟�?�BWmz������ 
(W*|!k &&'��ԈaV�8Jy�3���r)\e�O�$�cr�7�Q�"$1f|�����F;�^��31�J�p�.}PkLv�z�����t�oC�j�V�|��r�t>�kdpv�jb���g�d�m�}��t���v{���1u��DĔ��X`��2�QF� ���!�*y��Ba�m�漆2M5E���6Z��(c趉E'��/�)3���;��8��r|��]NL�{�Ag��s�_E�����e8Ĝ��&�u���فG��gNK�{d�{L�������Vv|�q����wۭػ�nY��	�^�&I��ส�ɽ�ѩtf�����,�E>�eTW7�Cfj�KIC �����L5�gX�,��T��ǩ��ZGU2I�ʽ���_虼�ן��[�<,�k�����N��>x � ��;���-����t��ط�7�C�]�Qo��5���4C����Z�םFei�����R4�rﶈ��)J��fr�D��&9x�9=�[��r�;�@����Mr������+�������7���	9��G����ò�U2�������b���.LQ.*�>g����gO��	��XZ@��=��%q���آG�1�F\�O�L�ᐴ�Yj��R�bjfG���t���U��C�#��u�C)"�p�8G���ѐ8�	;��0Ԟ��W��W�9� ;f�_�^A�D/��*BJ9��"-�P��v��Keg��P�`/�RA(&��DP�e���ʈC!5���&����
�i���4�m y�4�����dF�d윣'$�¹��j9�j�)�� ��u%�v������4�lO_��!�*]9��-������� q���������i���?֗�
�U������c�RKV/3���?b5k��D�v��І��c��M1:�"�.��qF1��o�-C4���M ��a�E�ꃰ�۞zk#��C�,/k��(�o�g�:MVE=��i>�OugТyӵ	�z��XR|�����B�y)Y4�M@%�s&L���XR��������ZA�uZ�I��"�g���=��
l1��V��?1��t�eW�͵����/�S5�6�b���t�zaC;������	k�Ӝ�;pq����6%��1q��A�)J�.��ly��6he8R�����5Vi۽Ny~���C:v���G}� ln[)�ib�����k n�quV���X�����cB�JJA��:nĭ,B����W�'Ck?J�6
��|OA� y���{	t�  �����|�r�
��fn�Z��v㕹n�<,�Ȱp�K*��**�9���b0s.k�����x�!]��C~�NY�E�-RKnE�|���7���pX4�EZZ<#��K�b���"���ݲ��>J���0���(�,}y�@����q�ta4�5ґL�!b�c	��J��Ճ�$ӂ�t)C^{���5�*��&��,�&�bP�afx{��uўP/6u�#�_�5�8��t���l�@]9��]3���U�|u�12�R�1dw5C�a�h����no,����JK���w�w�����2���z��P�|vK����[ i��<�a{�}"��Jq~evy�X�w�L�)�s*y�J���N�?��:V�O���]�_�D�$��F�#�Z��fa�MvaU�gz�p��5��
����Q���˵�,���*U�(��-��_��yɡ��T����� ��N�0�z !A}cnh{��,�R������r�jl������n/M5��>��jU�-wxX�vW&�t����[O�V�cpAY���sZI8	+|'Ђ�mZ�2���MBvo��5�(�y9��8�,o�#x�ϛ���^�C��(���<bڅ2Z!/����[\�A���"��F�SH�8@,/h-*�A!��5U���;����bFѯ"c��?��(����#��i�d��K����΂�q��,�n���,q�ROnrJU�!h�y�L�P�'.Z��Z���}pr�����۳���������l��-S�i6:�`���^�{��>l�&ieM (0ӹ1hy�Q Ϡ�}�@�?������ �b�F���Ȍ�b}����P�b����3�=��Z�2�:d$=���ѧI��XR��x�G��-��ٵ�i��2|p�+EA��	�K�DnB�RV]|��I��D��M�����NcF\n"�n+��5*���U��<�E+I��G��=�s���"�e��pe��3�����[B�4qV���Z���ɋiX�7�V����L7t��b�y��%�⎸M�Q�,x�~�ј��`��9M�ך�r���F��#�77`ʛ�m܉�͌�<y�m�����@���a�=Ne ��O3F��A�.-6*��rIz�w`�O'><��-�D��x��	-q��E��*���
�~1����%��RO카��A��$ ����r���� h{B�c�MH.�����u󑊇2�U��f�p����2?r_W��͹�	I]'���,=�VIƍ�3��vl��.[�1R�ڟSU |�����D*�~���ߑE���=dh����[^{u��LaK�@�R���?�6��T3�4��nZI�cS0�=�5��,�E)���=�Ȃ��e�*-Kۺ�Ǳ�e���9�k �#U�;KL~��t������t�NS�09J-��b&Xn�7�Q�7s�u>��Ϥ��U&�t�~��E�Bw�dv*�x�o�?���/�W�x��P%�	yq�AT�m*�z���7���Z���9�s])W���}����̂�Wy*s�I�D>���Ѻ㓺x��k��e��J4m���WZ_̉�ƈ��N;!?�Jq����@�f����s9�iM�̷��	{D�������Y��H��0���T��H�K\܊%��uR7߈ۘ�g�#)���!�t ۔P�W*�H(Q�B	�;������s!&�g�GtJ����,�m��X������Nt�J�K"NΧ�6��y�^o�/^��H~���ػ�o^S��k��uD�Y(��?@�s�ZN�D��������/0��0C�.��~���T����h����l .�dxv�lX�Vt�X:�,�6�A��ޕ���3�j��ߌ���+�l;P�yj��K`y(U.�%2��:U��Z�/�t
��3��*D�$�Ļk�!;����o�ɻbB��ه����m��G���rjp_� ���h�`�^�̮ԧ$ؕ��}j\F��R/(�	<��T�sn'������ǜ�5���X�\Y�@x����F+��+����U�N1n0�5��3$zg	�0�p�P.A&fvu��\���i�����G?�S}V��T0`S7����o�?'H�A�8�4�`B�`�\��M� Wl����3;����L%BL�Y ̨�w�I	��`,qx�'�f�+F�qVHsJ�;���;^��obg߁�;�%.��V#{�YS�1p�ڜt�9��E�Ƌ�>)`Lz��U�ș��O����<2��t�(�~W�>(J�φr�8s��e�S��_����(��O3�u�y�DTr��	�S�(���Q����c��+����F2:�72e�Э���_������A��X�,l��3�!S)���ə���~$7$�7�֥O�w�g��	v�Vg�$*C;��5���h ��A�P�6�jO�Hׯ}�M:����m��,_d�ۅ7�r7�_8m�(|�����Fd���È�0�?V?���W����P�Sd�j4Ѻb����{���D%����H@)��C��k�h�X����~޺�kCa�"�{}�6����G�i,��~�����6��ÿ��=!��4�������#.:֮�93�zs-㓨�A8��N�C�ȵt����W��Q�")�\��z�K���Q���7���<���׋���FR�m�S�9u��)p�	B>�EDb����m�U3��<�`��C�3���u��i\�~�8�\\���<+o����թ���B�#�&���Eqr6�6t8a���j$88w.M~W}��?Ԋ%�N�� H��L���9�v;���t�L<%ۣT^�2�&��W�*3|�2�x�ഽ���u��P�����>�f��$�GD��;���>��k�w��u��nB��F�FDkq�n�;I��^�����W�e����Ӌ��OQj�����^_��gp�������]?�&� zH�.�h����>Z�"ǅ;�y���F:y��ё�ku̅�ɺ=�>��1�۝�Y�)ǃz���)q��(h\�o�8�a7�:����e0���T�r�Q�XB�����f� �T�૩36O�L��0�R��iŉ�D�,7�Y#��C�Z�����%·�CW�C�>ޯ�^k��8ma���/��ڸ�iS���AZ/�ш@���t��Nͽ/����~���*�K�ﶾ�V���^kv?��#���W����qk�;��ѯ�,.�S�#J��4ғu�� {Qj3,�H�`TZ����Y)c�**4���M�c�����,: ��7R�����%Q�}3_Vork����MU�]�n3紁���7 .��煪����}��4���V]�����t�j�x��n�]�uFv��ORf-\�.|�bp�J4���t�9��/�P�����q?�:��-,U���G;�7% Q���?a��j��� �5�;a��ykV�k�{��z���;쯩�i&P������$�*P1.jӨ
��Ue��	io��e�_Y�[G�,Җ�K�*���8-;r��"9G�ţ~-�N1og=:���Е�,!Bo}c������ǃ��s�d�
}m.Ik��Lā����f�:�&�(�"�#/z���sv��*5�Q,~�,���+c�ieHH�_�i*�BjB=�/l�?����A��{a�!{�@���WH�@�1C�~v֙
t�b�SN7:�p4	������M �%[�a�5n�(s2�J�E	��<p�Ֆ�bp�:�ѕ���}�^�҆>i�<������,]�X���=��궿	��؃�kCtBY�z�>!G�j��{r^�[+�2��g�yAy�;E�/)Ȓ)���O[!7�JtG���C��+4�,z�^���쾄t �ds�X	5�oz8KIM��8[�抉ʐol�x ��@���>��B/�Q��z��%�� ��X�4�z��w�Yf�������H��"��]/�Ж��DG�SSD�W�ul�8��qGd��g�8p��%��x���b0^(�B$������fW?U � xㄗ�=ݥִͣ�(��=U��Zx&M;� k9W�dĞ��ѕ�O�%i�,iOߐܣ����K~TF��H-�>z�(,���P��b��%���:7�&�F�ǁt�Y�=p�����9�ʇM!������><�D��B��X6���Y�ȧJ�n�$Rn���Y@k|�G*�Vo��?�k�
��A��T��s ��9d����Q	)���ڕ������m��:���~����lݠ���ag���F���"UҔ�q��Y��z��Іo��I+���m�M���o��젉h�<�zv�u����nx��K�q@��K0���܀oc�+�4��o�syt��H8 �������p�)B9�*�`����%D?���"�U�ф�ԃ�8�1���ndZھ�S��l��(:��m\���H��R�q'�W��J#�%�	g�-�m5�'���h�u��p))��74�2�MT��tq�������_BZ���������П@; ojp�/ƶ ���s!4e\�Bn�xu7�"P���!"�����Yfz��������A�8�<���iv��A3�./��W���1Do������j�r�^揝y�{
[���)�{nG+��w�`�څ�;��Jn�o��7�^�.
"��ӸI����a�����.l��gZ�_�ۋ}�1�f�f�L)*������_��<����a��Kf��HʰH��.w����g!�N1�VR���S�g�hq��@��G0bsgC�ei��K#ne]�� ��Q�"��1�����epj�旈�蕴%T�xUp��@�^7PP�����I	!0�X��gG�?q�f,����}�<=�E��Tb�jR��ɼ��۞���d�{9F^��lqG��E�|��u�����/���\Q9?K	�[�w�m��.�1��G`��L���4����DV8$��k�r�r��Z$�s������?������E�F0
��O�� ��v�;r �[*`�a���z߇_G��I]G�Gi�G{g��;�01��a�Pf���5u��j����ک["L����������	�yf�ULm�',��(k����1��5�ޫ}݌�T6�V��$@�;�B�k���q�j��}D���i�����HZ����嵀�Fj�"��d�|fV_��-�2���B,�6�h5��k@0L��[7����׌a�T4�w��kYY���q���Px���iNz4���vI�N9�0H���Ӻ�`�asy&�S�D6yBt0!S)��H�ڃILu��f���.��$�J�iW�K��u>��|�RcWcȐkw�(4�-����J�T��_f�툭�ty�J^�4���O\J��z����9��A�3����8`�U�����o���e��5��K�`";�(X�����6#�-�n[7؊ a��8yOMY.�\�l�6ӌ�x֏M�||�"�|��yVJUQ��'>��HE7�	ʚ`=K����8�8ժ�`8_������Ѣ��bo�<�g�WE�Or��������c$�I0�!A`�2���Ƭ��u��|Ϭl�ή$�x*Ғ��!lX�Hk��i�� �'��{`|��D�����Q��]
'�:�GE�ժ�3����sV=��J�Vįr �9� ���l�`34.,�K�P����P��~�Q�|V�E�I3{ 3g�Q������vH��V_o���M���/�4�W���P�R/�����0��c�SG��u]/�	,�n))_�Y��[7u�{X�����#J�t��癯g8>��^�1w�/�<�b"������Rd�%$��q�1�_L��Rh�N����z�/h#J�/��fH�`���,Vd䔘%��@A�"0U�{KLp:=$�VKC�6�@>�^֛0�,�N��>��A�5w#<���޴���C;,���d��7b8�ϒ@+⬅Ņ�6H�i}8����9ٰ_a��7���ص �7 Rs�D���N%��1�p��lCsd��DN�u�{,�ұk�%tx'2x�BY��q��b$� �hz�� 	N�ʺ��2x��)1�
��O�'"�����&s�y	����yn�6ᘠ͞'�Ep�8���pݔ�i��.������2�GU#�1�mޕ�W�^QV�)��=���H�M4���̷d��J�]p��� *�1������{RBhc���������P�" �C����̲d}o���r3^�(bs��MyP�}�w~�\�A=&�ޘDC*���&|��}|$��MpY^NgË�C��q�@PR	�@��`�M�(�0�p��s�ϵ�A����8��G-�2=[&]�GQb�n��UJ`Z��(m���c=}u�^/��&�1�$q�O}2�5E����$��_O�1�deЖB.1�_~�}_�x�P�U��쳏����7�{M�4��Ȟ:z?�#ھ�`����l'�}8�����r�kc`}�8��'|�n</6����xb.��h�����EIr�_(�{3^�|?t-�8F
��
]]uE�� 4`���[ਗ਼�=0��]r�:O���KW�CY����	�/�0�#!�Q:��F�@,�N�T�������T��OA�������7L�_��J\-��+���xn��a��:/<ȒE�a�3����	3�]�-�������f�_Y��t���!���n3u�p-¹旸m]�oF�8j�q���ʋ-������LΏ��樕7�u7�i?8��}eP��j���)\��B *�Xq�=n�Z���ېI����l��zJ�d�N�h��R�?�<�������/��7��Fy?�KZ�U�Yd2��R_�*��A�àIC�Hg�� �>��t9�X��Lt��s�-���iΰ���s��]ac���HB�9_DR����4��|���i9li���ݸԶ�խx{���ӏ��MTY�EXGy���_ �^�.�@��!f��ZI�Z&��@[QЬKn�Rˮ�
,�08��&_��8��4w�I�Hx q�OU��[�$n���^³�C��D�|M�)� *X��L���w�Btm�J���x�q��[������mӼ��XFr�έۦ ����6���X���C��`)�C���5	�݈߂TN�u�N2�!��K*ws5�>��OL8leu��Mw���?�\�:�:����_e�!�:Z8�$���a��{bX,tK�pa�~pf��V�9"0gcLs�}tɟ��B��m<Rg�J����|8���f�۫1�%��J��4XJͧHL�(�Ұz�����Rg�+(L���y�us��(f�ǭ�`ɗ
O�q�R�g~SZ9�P�x��q��&~.$W5IC��`:��Ӽ�r����zۼ�$��SL�jR&ۭ� ���.�����}"ʏ3���=�^��
]�	5,Yp�R�!VC`�	_�a�917Ϧ�h���cau�ՑQp^ˏ�>����k`�%WPPW�(��w�'j��i��� �p��iX��"(&b�Wp�d0���_��_~�K�S��0@��-�'�2�#�,�1���֓j�{���[�m6!,��n�87����^4��hV�jC\�����~�Ωa�ڍ�<�F�l�$���aE�+V���D������z�X�����f��n.�'�u-|�G$�x�=/VЌHr�r�'9�Q�3�=��)�V�����1�����J��#糧��$����=����I�i8�vZd���B��3| ���W���Y��8�Ѥ@Ӹ�?)��65);��|pWg(8�@$��I1o�Q�����*�1�)Oє��!��I"-Y�k:b�F�t����9}b��M>A⼼��� ?�߭��T�py����rmx���c�a�Ma("F����Bz��I:�Y~����&B
�1����d\9�A9kWQ���в��p�4P^{z{�p�e���J��&��b�G\-� sm��"�Ջ�U�!6��ㄦ���Wh��I٠�Ә������AH������#'񀇵�c�ÙY�C4�,����W�=��>0#�YݡM��[����}�(|��hN�&)�(ɕ�&Zd0�TX&���d=q:��� x@	�\���4�STH�C��]��,� �`�&p�_RqhjxD�] yv�P<ݛ�[��[�*�&ެ.ҼS�9ֳ��`j���R�q_���Y��4�[��.bJ�u+҂Fs���R��|�t���{�.
���\�aD��9}2�F�!`�
�]ٷzsK��v����פ5�GI���W�".�)���!�^��G�e���.��B�A@�D`<F��lq��(�充�i��Af`6�$g�i�P�p:�*�Qb n�fӿ��C���e
���%� ��ݮ����;B)�r�tw��f`Bf��W�@�l�_�t����2��5���\9���և�s~��a��a@�aT�,*�N��Gg!<�����=�u�r��Vޢr�=�k0�ǘ/K�0�GYt]���g|��т���t�t��0�d\<��g�ԛ�#�"��gB�:��s؍: i��F���c�%��i���T6f:X�(�O���N�N�~����7L�,ãuHxLIcB�zrk��p'iT������x���n2xFƷ}�Ty�C�_��ü�Y!�؃�ٓ`��׃MƩ޼m����W����h���PPN�GMd�ԫ�<y}����1��f-����צDc5�u~i ���kt1vbZX�#�D��]<�Udb���#����VPc��xґ|y�"�ʚ��+�z�%�[�]BR*�������Bnpu���k��6H.�Gu�қ��ӍI���%e>>=@ ]��;5�Y��&�W{P.TEJ��y�����Ox��]�1n̈́�����ýu����i�U�Ȣ�=�_���Ns�۔)�H���M�G�p���݅�`�|z�AG�I�˃7�vt�ȄA��ܿO���b���('I�4p�B�y�im#pf��C"}� ���&�^;ED6'ݧ���j}"0)}���.UٿA�� 8Z�k���K_I0Y�����^�������pN�>x�h���H֐P�.�-TZ��80)�6ֱ2��TѪ���S�p��7�0Hnr�%)�ݗ��Q�)�ϊ��F4���
7 i�c3dӷOS
����
4�2�8]Z1o�}��p4�݋�/�f�6ׅcl�nmDb���I;�7�D����o~���Z*���k���+��X�F�@�e�M�o7����Uɧ��s$�@��#���9m	��i��iJ+�N�(�c�d-g��?p�j�Ķ/�Y����|�u��\Y����/ìCϗ���fx.�8���[o�I��0�C�� B��V�T><G�6S@�H�S�&�7�R�@��x�g&��w�P�lK�w������>0E���cJi��2��l�&�t����Gq� !���m��t0!I�)=�f���pV=�<��f�&.��%�������@�2_R�ċ��T�O	K���\f����\JD~OgzP�ŏ��"�"�?RrR)U�� ��^έK���
��]������������Y*�JeG���sk����$o<�L��.�Mf^D�Vx�p�(�:s7T������~IMH'f�|����������(�d-��Ͻ�<x�,���Gz���N?���jE���O��d}�dd*��P�%�L�4�q��_�\�e��d�.ó���q�=��fn�'�g�P|B&�uf��%ԛ���j�:�������h�c�;n&��k�v���$����/-�e�;�����vaʢ
V%B���TZ�9 �t\�,��O�p`�jg��Ę�2�,��6>K5�j�^���^�;9r�ߪs�1uŤʉ���Ib�c���E��q�8�2��+��1dú5�8�t�٧!��6,?I-n���ʭ�ϸ3iz���c�j��I)Ga���Wo��J5~��}#o̺�iI�8��� �ve#*�n����mT�(}���K�(CM���B�6x���,���o��*�'��bRl'���;$�q�y��5���_��5������t6ֲ�{3I
8������xQINm��c�R�����<�6��cU-Z��y�m1���	�4����	fg%�[|�76S���г����8,F(ܐP֛�8����t�������{zm��������ye0r�a�n����hF�Ģ�B���R?~'Ct0>h��g�>"��#BƩ��s���Z��6Հ��T:��+���4&\�W��UI��(>���E�S'5+�ǡG��5U��%��{T�kxv4��CɾJۆ�B(��P�C��R�׊A����oO��{���:��x~ 0���oUyF���l���"��GT��D�e�a���d��}t�4ͭ�=�ȭ'��V��H@�m%AA�<������s[s�I;� ދ��{^<�(�Qe��ؾ=8U,D	%����A���>�	]tGR�aᨱE�p')�%�iO�v6땁�%�"�w���x�1���=s]:��]�A��W���sH�nQc�3t�Ք�*3�_�,��
�1��Е���xr�~��;1])���}����5�(
,�s�-5��<�,|�'\��F�<t��<���Xv;�W�e��B�r���i�������HP�y���U8Ź�v��~��D�����.°%�S�d��=ù`'Ӡv�U��㉢"7^�Cy�Z���aW�z�/ė`u7��w�sГ�+���aK��[�SGğ��5*�r�װ����D�,�FT� ��myb7|-�V�" ��D�[���y�i�!��Bb>���!� ��H__����F�=2�j��޼����5��g��ݥ�j^&'Xt�XD�D
qE:9y����hF~�'���Z�[����@Ƥ�y;��\��C����"%�$<l��8H[�\�X7����I"���
r<nE4�@�y�r�O�@`E��e�� ���������h����^U׳I��/D��n�Z8��Ts���f�D��}zy��(�x9�ILM�б4��&�\4�y�m��+�����p4�y�합�H�K)W�����֍�,F�;�kMv��3��%*&3��k�ۓ)!(�l��eߺ���9�K.X�����rxK�x���<&jhc����EXUr6��MQ!�jP���t��ޤ{E�h$>I���H5}0���-�}�)*�}�A�N{@F�b8��jz���2|���1h�wn����X�q��G7+��G���P�����C�Gze:��-a��}�$8U�֜z}��J�m������'��E��gn.WC�uK��ШF3�C{���/p7��ɥN�@��.�M'�0]/��ڏq�(�)��T2((%�)2�ts��P��Wy�0J�T���7��K���i]�}b�gg�&�z��|�8Bc6�u����Lqp���X�МJ���#\]w�P���6���¸J����e��%?h����N=�b�dd����8��-�L6�o4� i��(�xs���������gq�Կ��3q�[Q���2<lv��q��M�%Չ���c�kV�@����U>����+.q(/�T���+OY[wf�� ��S �qt=�{����5����ӌ0���0��T��&+Τæ����VL�k	vN8�Ȧ"3"�A>s�`���*����I�q�x�� ��尚� "ض�+�ք���\@��/,y���jL�B�윅U�S���#�s$ڢ�#�o0�"�FXZ=E�f r	D�L+����7��������=�� Հ~���c7/zd?.7:J(����:�u,�	F�Ju�ћ<�tH>�
��� kl��^(�>+���Q9�mf�q�>M�s����7mUd7�����c�X��7�W��@l=k��>z�O7�T`4�*��@��/m�$�ƨt�>���L��T2'�����&��r4�m��l�=?.�/͟�(4����Mİ�Q%O;�u�-����a����b��H00��\�:]�ζ�w������ğ
'��pт.��Gx��=�V-�_DQ�u\y�A�oNr�`�AC�}���|��^k�����-2Iu�5 /���BM�K����fk�RfՂ�H�u~�?�E��И�Q-���]�@��������16�JSV�o5E�������O��'��eP�c����֖WRK!Y`��6�ywIXZ��<�W�1ԹF�!g>�^�nf3 o�����]l_��@p��#Wsҷ=5!������BzJI�^j43��Ģ�3�I�Z1��{�2bʥB'*:���
�4U��Q�9��Q[}/�_Cj�R��^$"��2��L�_������������+�.SS�Z�;G��yO����`Ͱ���N��gz��5Y�;�s�͘*CH�Q�ȃ:�Q/�s�����x�ڿ��ɰº	%�P�=)�ܳ/�yI<���կpn���l�m:�pE{I&��B�=�Ԃ�$�E���EY��#�v#8N������ϗ�� ?�>;\�J���EF�栬�޷V\�+°�Zf�s��Ǟ�fD���:-7�Z�����f��tȁ,R�����MQB����y�'ĵ�]-�Ұ!Y6_�����7�����W�?0U�d�$�N�L )?uN?�^ߘ�).9�A�w���?���7��� G	<�~Sn�j���!��_�5^fVt ,� �+��i�&�}�	������/���"�G{V�Af�8�p��J���*�<���8K�84�a�c��QC DëO�����]��B�Ϡ�fق��q1������Z�o�:0�����gx}+�g���$�U�S�+���5���z=éմ�⭐��Z�����G�k��I����:�M��9N�Y{���JAA��ɼ ۉ0,��A��U���(m"��18ݫ��3��Oob�T�뢐� _a*qǻ*���~���(�m��`aCg����>*1�r�����,��dl����{������y�i����M,Q�Cٞ�U��P�l�s0�*wӨ���	ɐ���z�d�������T�ͥ�����޼��{������ NU>�#g�P20�sC�*������\:��W���m�OY_��-&����t����$�X$wC������9�sP,e��)��?���R��)�yb�N�\��ƔL>�6a=5qX�����=D��s�����C6�j=xAB0Ð�Kbj#�x�&�݂��v>����渡A;0��1q5>�ҳv���L�?&�Y�q�q��'�XhZ�Q� �J�INѼ�l��#�"Km�H��~������߉�IG�G��
�R�Gs��$�&�t|���NxЩt����/�7*�_)��-q��
[R�}^�����8�B��R��#䫨<���)Xe[_�����G�'[��.�ƅ>��EPxt~g��N+.B[��RT��n�Zŕ�*���N�&�g]���>%��q��I���a��#�d-u�,|3���PmպA��fF���d����+I�~��&7<��s����4Ty��m{�(g�/�(���\o���'r���.���A�Q4w�i�vNG��f,�N��	��v����,�ud_.�#?��n�����"	n~(SLJ� 5?v�h�}��Q?�P��ؗ:��^��a�<M�>-b,�����i��Y�Q8j�X�?����;/��?tm�%4�n�Zh\��8�|�/HǛMG(�a�Dtߡ�ʗU5�V$Z��R,�.�*3k�}7Y0�
�	MA��y�YA��B��>`�����Y�I&���%�?���?C�`����4
�A?��F��5��}�Tʗ@
�&oA���/���
@q+�2⪲p,�Fv
�Pq	F�͜m�/b;hj�i����;��d�"�ݐ ��p`�V����$U5���J�0��_9bZ���2~(��HF<l�y�zjH�K�1��o��3����R��w,P_=!A�n,$�=�/���z
�ΉH� �J !��^�2�ަ9������ލM��NJ���.{cYj�ƗS2]�%�4ے�8�tHN�\B �L�� �pq��xBۦRD���5�Qq����~4�]��zI\,�>\z�Nf�^�˥��u�e��]F����9&=l��$?��<p_L 9�N�FA�]D4���Β�츪,4w#�����-Xa�-�0CX�R(���೧y6�T��/�*^qkd]	QN��;�s���#����ì�X֌�����y5P���n��}���kz����8�g�MebA���L 0НO[i ?ٺee�z�z4_�d$�(�>{|�Rn�@J�F�g���ݦ��l��y
����꼃Z(&��N�0�ޛc��
���!�̉އ9�x��"�9�y���51��n_�}�S�{��U�bށ$���;f̦�5�ki��ip�i/,.��ܦep�~;3�P�r�<�p��F��J�ֱ�J�U��/��eε٭��s(75�����6/���'�0�r�|&?I5(�.(OU��h�;��	���t�;�Q4|���J�?���~���&|�?E1����L}f-o������ғ�ZP���A���3��?�EI���
M�gB�
>�T���#3iQGH��-��!)-�3�[Y��n���R�o>f����9�(�Ne�^wY�WB���d�� _��V��k���V���_з7��J�}*�~����#�PQ��d��%����
7wk�2�^7�ۃ�;�&!��|�&oj=4iJh�c1���Dj��C>�n�]�gz�g���U�nhx��P'!��c�^�_Җ	d�!�6�.�q�/]�wo�/�o#'b��kS��a|�{P���9�eIyc�c���vT{�Y0,��CZiN�\�d�{VWl�L^��?� ��ٶ�0ɕ�[X01�#ȺXc��-]��aqx�lP���/3U%���-�U=w�5L��Q�致�kj�	��R������k��Է�3_Ҕb�*~|��Ee�OPE���1T�	.��83�{]�	�3�#�7'u{�������aP�|Vk�ٸ\Pd"��mjm����8��G	��F�LPQn9Z�k��F�Nj+\�*�'uV��=|���p��������2	�i\�����f���Y�畜��e:��ƽ%d4�Ɉ��c��=�vE�Ǡq�f@S;�����3>��n����b���%��<Ev^���J��*�:�$)x5n2����)���M ��F^]l�a����	�q�d������Uy�V>�_�;��?�R�2��:��O�j���|t�`��~��ֺA�p �I�L�Y��X,g!n;9�\���{G��tF`��x�_`h�q���ݔ3u)6ԑ��-UƗ
3� Ө�y+��ޞ��^E̼���;��ެ%�>m�3����:�����O9A��<�FV��TYo�'�ӌ�2��A�����K8+]�1x0������9J�}q=�T�#Hg��zf�����R�Z}aX{Q[X�H [㻬ή}( Y7QLH�|#�;+�m6��W��T���.���n�E��j8���t8�o/�t.��!���!|<��'��Wr㪉?_�c8J�{�y���}:��0/��0���[y�s�9D�\��,�pJy�&�4�,0�p<�u3dXV�������?��q�yU�b���Q�׻в#�J�_x�����/8���y�r����S�믓���S��gx�3萭�XΧ"dTNly��e���R��΢�"�l.���C����4��h3y�y��Q�(.R�X��&�*���z��N���[��Q��Rk�r�`v6x�m��y
�|�'�r[>��/�R���������R�i�\���:K|�y��Q�����*L`ʛ� P�$}�s�;��1Evcƻ����$0���n����D!�P��/�����P���ԁ4�=���;D:[�yAG!O0 �ȡ<=AU��oo�G�{�;�=p̓s^ag�g��Y�W���fjVM��O:��z������f�?�G�Ij\^��_��GE��/�&,�줆˘v�����I��A(���w�n�4j���ˎ����T�'�=7�Za喙z
v%�Eo����ğg�r�?��;����;���	��!��pB+7O؁�.��ĩGpn`�	��.��TY\�T��?���^Up{a�
��f���jK1�~?��r�s o��Tv�c�%�^�G���j�U�*u�Ň=Z_K5�zT)y�H�yӠ�:�9�ù�����yF�6����g>�-�}Hv�(@?_�}d#���T�0����t°�����2�ܨ�I �Q5��TQvϘ�:�.����<����)֎��X��BY��=w^m�Јg����tj��)M�H���?Z�p�C\�_ �p�O1�SV�=��>J׎tx���D!����9c���u�_^'��Φ��xr��wHtLƴ9���f�ea��K�"bbj�i����g�l���������D>+x$=X	��ʡ��F�OfÐ�MLF�5��iPoF�V�5C64�8����������X` �;�����)٥�<�,��]-�	0�O(�
d�SOC ��V�a�"���®*�����Ryk
��Jl�Q��ֺ�%Q���Z�A�����(��!$���O kFd�+#�cN�GŻ+����ɋ[�l0�'bQ���b��^�_�P/�r[�C��㱥l��
j�tl�1}^p]��i|yZ����}/��ـp20���RYY�@�t��=�7��5,;1]��-H:z0��-!;�T���5��W8�K�ңL�|�$�����H���Q3L�P�]�@���/�� d�k�m�gWBǀNHm(���y���.S��^�e�=��\^�s����	%����m���39)�l�w*? �k�#�4���(���у�E��g8"~U�>dM,�D7����༝��Z7�����Èq�n�;�6N��a���鲼�:�d��PEk��w!]%Na ,���wJ�9�H��P=�U���ܟՎ��b�v��������yڳ�����H5k��0�&��GK�3IWg�"��c���U@k��*y��YM�?��X��h��_@�ժ� ����S�f^A?ɡ�Jd�z�t�����s�
�����n����KXyo�*�ݽ����
Fr�a��^٘�/�=�
51R����t�E-���sx�@�p:Kd�L��P�	�O�r\�#f�\��*	�c���rW�R�̈���ɺ;^���<3:������w�`�L�P�sڅ������}<�o�rte���vg�Ir�ɀ���+$ZզJ�X�G&���L�{��Y�;��d�����tG^5�1�K;b���;�R�e���"/-h����Ē�Sғ��+AX��|B��-��)>8��M_h�8���k)�!�[<2�[��~�W}jFj<6��@f�h:`��\գ��#/޴8�l��C�da��J�t6���c�"(�
�-T�.lm:9_7��/�� u��U��u�O����ZX�T��cи�tUVd���I�uZ�HKI���z���e�?ߺ�����ѽ�ЮJeS�i���
����]��=�k&a�6�F�cp;f�[L��\\�d����V�%%�׾jQkz1�����~��zx�����~d�4~3�)$
1�]���P���
��$,bٸ��6N�������gQ��D<��*����mF��NJ�2bF���Oy^T���Ϥ4�8�0����[�_�o���l{��@F���\Ll�3�N������������]�	��0��|+Ū2����$�X`F7���5 �8րwU,c��	�ʋ�)�X�7ݰ�F ��~�i��N3;|�P����O��r�Q.�[l����X��*����C,7`�!��Xpɚq����VR߹=$Q!X^��b���*׽�aPCc��×�RͰ���6�˱Z?FU�Mm���(J>7�Ǽ�I��G�|�2����U�0��`��u����Wh��Z�n�R�L��C�B������|�pC�n�x&����H΂ַ9�;'�8{����3�=�ݨJo�
�7��2�G�������|����^} ��f�V=��k�]�:r~�_���1t`�ze��6�G���}n�GI���/S�x|Ӽ�gX�k�I^�E��G�2`����=/eUOM�V��.�o!�%h���l�?2x0�=�=�N߲E$<M���xt,�1�z\��f����}�I�t���ў��dr��o���� D��X��+g �b� �]m�u��&� �Wղ��������2�nK|Pɗ���E/+^�	�C�8*�+ɲ&�/G�@��v������R"��Hd|�����p�E�~XhÏaZ>lu��
>l8Ǜ_�^K�m���ΰ]b>O�.f~W��nz�����OcԲ$m��H�X��h��b3D:�BL���Q;'����x�s���~�^t �g�ye#,�~`A8&Ά�@�+;y�vb��7G`�"6��8n��dO���.���c�� ��s'E1��K��{qkе���	.j��%CK>�f��$�C�?��B���=�2��]%
��.Ʌ��PO*ťa��Y(5?�lh'>���
�L�4 ���XK��#�F���,��#���3��s�#���6���^�*�%���uƮ7���;�ݞO9ù�i��E�G͞�cF 72�y��+B�%ry5�Z��Ж�{�jh���H ��J{�[��9�pD������鈁������^��d��h#�T���]�7W����������+����7��V���I�x`����kr�u�������y�������]4����U���+m�D����R1��j�S���&+��6W���}ϩڞ�y�i�<�h��;x�3�U�Ml!ٷ�j9��q<��Z�Eqo�N�<��=�P8�j�o�KQ������%�'oc���i�DD�K[=���~����#q��&z�uL ]|���c3�j}�4�G�Ey�L�@��=�K� �۰�`��t�d�?�N=����t`�-��4]O+xz>ř��'Oy��-�����ر�s����*i�,	7(�&`;c�#�rˮ~�:&ݬ�EI$U#��
�G�2&�I1�R࿰,*9=�Mi:�#���^ c�VXp/�}��g F!k&��h������,����2�;����u���t�ޕ���5M/����Em+s�`� �qa�X����j}���3�1�g���N��	�ݗAɴ���a�i����:k���k<`��?s�Z��ǫ9��J��t�����8Dy�NR���v:���mb����y�pQ�f���f�C��)���kæ�H�d�3�����qwf�rK�c	���Z*,!����)��8#��\�98�n�_(���94���ղ���	��rV3��c2��&�0g%�4y�\<��@�
�ʉ��}_j����̢��=i�&u�4�~��&�!������C��<��s"�%}��2 !��m��صP{6�Ԇq;�d�!��"�(\�B�mۗ,�͞�wʢAz�."�~��O�
Ţ)OsNiB��B�/���P�o>e3
 }�+�� Z&�fu��VG���S�V�ˢl�I{6�5��)%8����ۅG'.Q�pn�sQ��K�*���t;��X�-[MW9�\������"��м�j��F \&1C��WG��JE�߀Bج�
k}�����F���Am�=~�}[P���� _B	����!vٖ����1uD�4`>"��e�R *���j)��!>G&!�>ʼ��dZ}ˌ��H�`of�ip>,=ӑ�>7�D�{�N>�-wt���U2�c�~!�B.7n~YYgߨ�6������L�̀t��r��"3�=~�����T�&'R�#>�n�A���� ��d���1@((����m$M�]�vY�f�r�$����L;�[E��P��&�F��8uA!݂����[*����#!�@Z,���nr����:��0�Z�ǊTC�<=�Q���n�{��+L�J³�>��K�(��Oe��hΪ���&Q�1y�,���,=r��c��CE����=�ˉS���>����(�����	ܼ��4�2��oc:�M#/2"8����Yf�?_���@D�GF���j=d����ˎH���-?��3cs��8�}O����Q��5A �]�>�e�e��$�˰�-����}�&�N���� �G��}V�,���Q_�����J[N�35�%��P��Y,���[ +�8n���:>,��j��+�Q�(d��P��@AM�-��Ew��ŋzU���SF�8��5* ]}����I"����JD�Pa��D�s�ԉV��D���k�I�܉bD7\�C7 �%�0|C��H��ɽez���RU�F���ޮq�~Tl�g�T���GJs���S^}�+_U��s�<�P"�E�1FD�DÃJM��{��N�\�������-�8��;Wj\����U0�Wسz؞�>7��^��u���Z'"z�n¼�as5�K��-І�|�te}��܁�*����=_U���ҍZ�q�#��"2۪�]_���TƝ���،]> �&�y���!��T܈����eI(��9���U����)�ݩ����D��/�m�VX��zě�����LU)��욇(���5H�#z�C.X>�4+��Q�m�[m�j��](��H���<�
���B�c�Zm�.A���;`��p*p�����F��x<qC���#��}����I|VI���aRVSIM��4����|��/�]�d�}���kg�����-��	�LQϵ�5Hm�-F��n�7�]^�WY:C�ć�V��A#}�I�[�i:k9�8�������>_�G)Q�I,T�c���D��G;�J�[z�Q�R�q�>���z~�����;�O����
�(և�~�# �x�����TЋ�o�6�+[�R]h)+\��Pw�LS�t�x�+Q���\j�lI���B3����lIdU޴���3h�E����C�+a���"j��]���	Sp������w��q]kz���J�"�W �H��|(ؾƛ�\YZCj6�QY;�C�A�=a���-�� �AVȖ��,�� aSF��!c$&	[�� ��D2���@��r��K-U��[�%e���h��};M�UTM��y�$�p��*��	���Ӭ�pZ`�G��wd�=d�n6˕J���>DYc�����@4��|��bK=��48��	[��6��h���RC�B�i%��r;Hq��E 8������yY}9�6����D�󰦌B�j�d^c��"߭��6� ��5H�:���@��\Y�[f�Z:��a����X#&����:&08Ӄf���P�J�4�s��>�/�w�Xu8{����{�!�fC���Ԓ*sʴ���,�3e���3�x�ܦ�(�NWC
Z�"�3oo���DWO�j�Q�1%jTF8��==V�������z��(����)S�������H����[@��v���^����}s���D*:~�R$ j����{�xڶ⬑:��wx��뽖�Y3U��c��5�c=��k�7�����Ov'׿㠔�t��m�xi�rm�R%��b�ԑ���-_��[,������� ��Y
^���gT$I���[/�_XI��6�c��	���a� ږB��?��3�����k�U��u����P���q��S�J��|�mf��
w�K���YGƥ<����'֐ϸ��FEX���S�&�PY�nD�a�qpm���`�F�,�ϸ,�&2	�Y�fo)�7z�i2��&Cv�m03�^��!�6}]�}d���(���o�4xD�|O���?�T��H�f�%�I9E1� \�R�'��_�7��8H�;���M�g�kK;f�/�PC� R(q��j���F��"ȶ�v��kH��ϛxf���єR毳�􂃟Q�H�Q~xhE6�'Mk���D����]nK����%"V2F��^_]/6v�U&���8���,.x��"��	]R�z�t�x\��+ER��I�e�x��c�����'S��ݺJ�nj�x,>fo�g�&_0\�򍻮�8�gj��pl��d�����w��jk�)�uv.}8�Z>����	w�O��$���|b����|�X���ɓ�����QD�L�^f�ʄΩ;4�������+��DrB�}���g��{�RN�}��!VJe�
��@�	R�@��t>=�|#����k��5[�0[�}�R�3h��J�,�'t	��H�'#��?�W6+��3A�����U&�`V�	Wѯ(���Mv�{Q�P�"��x�mDj(��>ʸ �$[C��4��e�c.�)��L��	i�k4X"j�f4@DFjS��T�L�I�����y������+𷀰��.x����+?���[/j�j�^3<6Uǲ�����d8���y׼H%��E����Q�����u��"�k�k=ӣkͥ'����A� �҃��0znv�Z�6�:m���әϜۭ� ���0�����Oπ���
3n�����r�m���0�7�<�ܗ�v>���3b���"@���x,M��!��}�\��x��KZ�HJ���0|���鵣~u+�׮&�C�� 9>B������տ�)�oœ�q5��9���_�����n�5k`S#ռ�i�7�l������/�wA���ѵ���l9���)A|�.�+ǩxn����B�>[��!�|��a	��O�Ը�XC��%�$~N�VP�W��t���ɺ6�b�����3�~��i��]�Ѻ�/�$l亮���)����i�d�d��֏�����X����ˀᆔtn�����t�	+�uG�bʏ�)%���/�v��}:"����L9�*vXJ��/� 񢗡�6��V��c�v�UJ@x�J��ܢ<��qg�_��*�� ^�p������銨"��{���A�,zӈs���7;��.�N<1�TZ�@NW�oLo��ѧ3�B!��<4W�O&������~�Ǎ&d�mR%-�^*�D�o�Ժ�B�]�o�b�����7�ԗ`l���>�"��1�!]䪖���h�r4��%�R��Q"�ݟ:0���=ff*������I�+)����a�Gd�Xm����D�.�A�ch*V�3y����l��Z���fhzJY�)��)j��a�-L���D�!$����C��2&X��B�C���lDKm�&5\n�i�~|�)tm 1�7���@?���J ���'�C���a�5n�|"�|�[z;��������xK0t�sb�U ��>%�l�7���v�>�N8�]L�&6s,4.��4w�V:I�)����1��e�Ꜯ�DM��iɹ�6t0�hL8hA#�9�^
�Q����xO������Yo�`���k����f.�
b;�
�0�nE4Z5�L�O�US�ʄ��6����X���#�^���P�}\Ѵ%,�"v���t�/P����5�Ir��[���U�bH��Mø���E�ru񅠠�W���\��o�[,��w���D]���p��ݺ�p})���eD�Q�!��8٫F�E$�x4��*�EV�5�"x�P���eEB��J�U�/�Y��&��R���?�:Y��Mqx/a<� ��k����,�k�_0u^<�S��Ū�},��~u����77d�+�X���!�(3��ƞ���%]G4EP��W�g�FCm,�h�H�l��:IЪ����	��`��YH�w� �-ٽ�m�U[Z�	�L7������y���CN��܋������ᘷG����\�����Wӂ�]�ԟԄ���IJ�J;�%t?iѓJx:�p�1oK(B���˜0��5S���; H3�T���H#���z^xC��9�,�B�0mb�����K̈�G�E�0�wOM!1�W4El����#�Ҽ$��:���ll����V��������G��b������s🈌*���8�*�Nm�&oq3��'�J���PX4mˋ&Yz�^����y��.�.gڢ�2�!�/9%���1I�,f��-�i��ƀ���7��+Ҁ8)<�e��L����ZS��M�q��п���E�.$���ث�� ��<�>1Nr�t���{D��̒D�~�^�:n<� �B`ߎ��d������FfQ`��_�D�!_�pQ�J@M�7.a�b�;�֭πb��W�������&�'؇��I��m��тdM��)C�jם)2�G�γf��&]��j���$�$���|���L�)��7�Z�?xV�����O��
��x�RS0H�J;
�:W'�mߣ&�Mc���B e�x~��v�Ҟp�D��x���΀_P��bYvh1�z�5$�tg{:Ш�v�?1{*�y᭎u���`a�i��8���y�U	G ��jj�s�hZ*9@�88н�8=%�Co%:�p!��MH5���;0�^MF6�y�q�ѷ	��W v��5���(Bs��d&�!�@��ke:�z~��Җ���(���k��c L:�Z3QB����^�	sh�9�����$}�ٲ��>gD�"v"DKǿ����	��CCH;ص�}M�p�tYzE����Z���|x)�D��W>�L��zx@��V�gT�@"3�S����/��fN+��̙|H�h�+c�%R�ٴ���W_x�� ���P� ������v������?�NӁ�����
C��ȫ_kx����~
�B=]�aӨ���J�Ge�5h>��t�YRm~�:�W�1[D@�c9���R�/�Ey�Y\Õ���&=�Dg���*��~1RdBf�x��7���W��P*�V<�����U2�یh^UN�����k9�����?�n�D[P�R�1�828,yXY���A-�Kk|e����-6xe�/.��'���<���(�DP욏<���jT��g�õI��0�t1k���F�¤y���ϲ���B|c�_��ν#MW�%2z��_��ݗQ�2��mGv���>;W2)���C���i�t���Nz���9Q��P�2�u��.��¤ʛ��FL
qޢ7p;��\La�uy��wԝv��b���d=� tҩ�k7!"���Sa���uO�su`w,as��!�v��6����������p2y��#�!��0T�k��m6d�W��Z�z�E��L�M�u��րX��>7\D��xZ��R�]���ڜ"  ����Ǉ;�z���� �� ��Y5��2���17�r{yP��cI����W�Gş��ǔ�4��+3�z���q�if'�܋����b�pqq�\~?���E����vi��!ߗ+��
��'�hLy��:�8*T�e��U`���Z� �6}�����<�
�k���>����v端�z�wp�`�_�3����5/1]�&�Q�%yT%s�#�)�Z�a�󭗕��d�|ͽ���wɺ�k�GP���	���t\�&'�E1�٨��	����|��抜�H��'^�rz��'�Ghr�2�wb��/���pO�9̧ܙ���]�uT�Ӟ�P<0�=�X䶲���)֌d_Xb�*޽hA�U1	��҂?���TԐ�#����9��H?<�xС��`�V��U�6X8�Ś/h����uRG�u��h!c�Q,�I���B!H4nou%[�����O'@J^>y@3n�}�NTrp�>""ߥ۬m�=y�=HV�P�"|�6_�ּ�)[X�!p2�K�����o�W��PN�K%$~ +n恋 Q�]Vڟ�&lR8R�O�w������kq��p�ޘ��7����������Z��-(1�1��'-���F������vΆѺ���l���!_X�T5���:�ӵ�(��,LS�n���"��(�����>v�ҽ�]���WبSk٬٠���g6��� +��c6�_TR�A�A���	���%�;�=�R�>i�w}�&�K9�v�n��ɸ~Wm��U��~s;�G�Z���u�2���=q���vj�� ��Pݠ�C0ǌ��Ix�ϯlI��+��B��UO����9�X���aV���p��X��޿|����
ѹt,�PDf�w+$a\p��n�,�{*�Z3��H&܄�=����0Q<���'i�S�W���b[�,�o%�=ye�x�d�v謾gRy��e��h��u>��ό[��j.EMJ��C���c���I�B�ٶ�^ϋ�]U���f���xf�M�����"�%rd�O�
m���c(g����l�@�d��o9��(�f�h�|�V��I����w�Ӕ���'8���>��Avh�,<�"veD����C
Norē �4�>�����e���+�J�\�8������7����Dz��h��
��<����>S�bL�����u)l �#N-w�$�ѯ�k��"��:=[% ߐ��?�XK��/l�7{Ş�Tq���yQ3aP;k��jەm�8%�>|�� `�6�1�yg��0�}+�OB�1��/E��W�Z�;����1��ɐU��<�z/6�ri��f��t��X2�W?�&��lW��$��t��jǏY�ׄ���@�ȴ0�����r9�M�U��5�'� "d��Dk
��U��L���%�{D�T������5D����_�d��H��ϐ�\ �ւ�Rd��V�r�餷+?�CA�vl����1�<���˔1�RZ\m�xw���R ����I����]�g����}��u��&+�@$1�ڇ���g���ƈ���@n �Q�$�涆F����W<{�{�
�e�%#l|�_���$1��W���<���s���������>�P?c��N�p4ο=W��wdo�Z�ajҀ.��o�DP�c/���x9U2ь3�B^,��F:�c�k�ڗ\jBz5��N��đ�����)?A'��|������H+�Ҷ��S��= �����}z֮`�4c񱉞�h�t���?-��^!�opt0�ݳ��N�~�#
f
�aUrA����}G_TK��'d������{ɕ6�S g�SF%zF�;3�})����m�7��`ʙ�d�/WBi��W�O� ���\�%�A+^�te�7���2�R�P����M����o4��� �t��lJ_n���b�� [�R���? `��W��������g�ЯM,*$V>-��4W���Ib��o��ٓi��-1�2L$VZM�Ӝ#���M3�]�o��
��A�vZe�3�g�����o�[qɯ�[~�H�#�a\�1��x�ӭy�5
�� �,ਸ਼��$h�Wl6]`���]�w$fc��M��
Es�H�p�)���ډ�;@��(�<��rn�S�΢��ȱ�u�>�k�/���v	`����~:#�r����vp����C�鰅�и���{�U,�N��[�r�>b�G��%l�.FfU~&(�/���Ny}$XW$�~
����L��ۼxQ�`��8�P}�s�Ջ��P�32��+�k9-m��/d	̗cУ�K��lɺ������
̵2y,_���Ui�w{·G:g�d	 v�-ύ�d�q
'�+���jO���Q����B9SrM��������7'b�O�'"�����L�b��q�쨢�e���S�G�.�\;����y��4P�]��`��N��^�Ά�6P�9n�r�5#�y[UI�*l����^��b5���R�Osw���'��EY�i�{�/�2��I�|}Y��r+;;	�8�,S�����8}��ڴ�Waf:t�9�c��� ���~Ӧ���y�x*]����|��$+~�
UO����9��DV)w��K"���N�0�xJ*��xK��bs�nz�h-V%Κ��8KD���,�B�@EX��U�f~��p���">���z۠V	��ۆ|��-D��]��[`i���d����ɎԺ8.�7߻��Q��:�eEC)��%�������3�6�d�l�W��̉0Xȳ��U[�5E�\'ۧ����b�ic�)�Gg�r�@ǾX
mz�e�<�p�J�-b\��<C�q��e���H����`�W���-P	R[�a��{'�PS�
�T*kޔf�@��K$mߍ��T\���<�@+%Q���̼�F}~}u���k����`�o��T��Ҵ	~UscBXnJ��;��V
����"z'�VzI���Y�5M ����E�/Nv ���J�FkZ4.�%�w�k��*`���L:�b!�2k�U��+#��Pk�=Uӆ�5��=N�j���$Ǜ���5��;i�ySV��H�iz�z(:�S�o_��Nni�N�)���c�j�A�|'|�� r:���H�Q1���	n���y�J�V��Ԥ����K�F7CTd�]?��*#}������HP/�2�c��f1L��kc��Y7�;�O�c��ן\�;L�$�#��	��R�u���ɧ�[;�����k�O+��'m�����Ob�B��l(�5����c���'�<��p{#Z[�v~3�I�%u���q�8�w. �	�ҲF��F˅��	[��X������v�����$��g�j����L�t���s�����YCpx��EVJW'�5�(OّH\i��Tq5�cŀ��*x[�R���_;���/��6QQ<�X��R/g����+��6�1��~{�n��#�߂���fY�C���v�6\�A4�������\�뚞R~h[�����~�1��\��4���{:M��W,�	��F�a�*��Z���,08�[�Mf.�E1��,S�l�D{�� �:�̡���.�� 5u5���浕L�����I|�I5¢ib��(�H7&Y
�{��X # (��cT`c��O��
d|��Fo+� ��T��+}����-�_[��b<�h�[�CW������t;K;9���C\E�����c�<�b��ٞ, 1#Pm�;o�1
�"���*�C�@���	V���&�N�� �	�x�P�6`�M��V���d,"C[�ͯB�ن�$��>����,�_�#5X�.���vyʃP��.���xu�HX�c���7�3���	�~�V�H�FbZ$�.�c�1��Pu��
E[��� ���D�@8:����9=a��TҸL�m5�W�iD������D[��]�ŕc��ѱ�����^tӤL#����M.��e��`M�h��fT�6Et,�J���K�9I�&��l��w��?�9\�>�56>�y�h^=n������^�<=����7#�7}?�r��XK�^�v6Rz�"Zum�-B���8��2V8���ב�$���WY[�S躄Æ��2� f+N|�Ɣ��m{3��6�r��s���2X]�7�Ĩ8�w�zj(��>�Q�}lp��{/�B�]LrO�,w�;b�ؔ��e5�{�e�w��B�qzi��J.,7�.���r2��X��$1�Mp�j'Em��"K ���'8!x��<�_Q>�)�����ŴP���Oِ�H�ظ>PV72�3��� �@��_�:��{B�A!�?|���q�n����'�cЋIW$B�
?��2���V��.�dNX���
j��-g�'꾘H��E�/w�C�b��7D��[�LH�K[l7w�a$L�:����k��e[wc�JmzNM��#�
���M�9�����p\�l�:��Ïk��ΰ����2�^�Jf�2Ϧo;��,��:��j�#��>P���i���h*آ;�o*+�B�H��`?��;Ek����
㢼ړ�мƶ��Հ�ة��S�9�R.��g,����M���!�y:^K���f�� �b�(�Qm�P��K|��(j�Ta�!��!�oS�װ�y���4�$.��z-Ј17?&`��w��B�2��,��n�g:xsh�d=��#[��y]���!&���<1�9I����,D>S����n��q6'q�3�L�iuW*8-��l�n�@p��wfW`F`�xh8T%!t��_��{��9���4�Z��r��O�ф��et�h̏�9t�F6�!"X	�x�.�HL��֑��f�?��a���X1[Q��
"�A�NO�  ������I�eK9t�56�"W]�8��ƂG�b'��,g�e���h��l�����t�����֌��/�#W@%�%�&F5ʙ�0w�4��KD����i�"�9������çd�����ز��)�2fI�R��ر��f����W~�����Bg�q�>���=W����p�]2s���1��>��)<�!���`�Z�^$���[k�S�	�A��{�@x�>�i�?A?��5s�Q�{$y��a�C]�� �;�y�ugx�1����<  ǯb߾,�?�w���Ӭ�2���S+L���w1dl�,����'�Վq�����a�e��Gt��D�&m:6���W��!v"$�;M�l�d�G+�j��q/\�Ͽ�ܒ�"\􁅂'��=�r���v���T�R��ePA�_���4���.
�XϜu�O?������*r������)�ەm���2$�3o�迭��w�b�	�R꿺��"����vFP���3�҅�j��9S��-�f�b	�1OK	���L���侾�s��S���Cٴ��P�kba�!';ǎ+�գn�'�]��t�|��V��ع���ʠ���(a}����)ʶ�����0�/�o��'=�,n ���-��	�S�_6N)y�Q�.�F�	2��o[y���'J�̨ݩ�j�"X4�C�K�G_Q{:8�B�㑆,3y���UDj��bn�b�t�J������gF���V�"_�2	;*x��ֽҎ���Q��Jpc�/f��d2�~�[5��?�y�yO9V�7��j�0�<<̴�"2-?��y8���힂̐���t�ݚ ��O��C%k�̫����W⌕P�B�l����΂=��P�HL�ar�;tϦ����D�
8�׏�و�R�.�q;@�{eV���@���c�n���&�2������9��^2A�����^JoK��?���>��'���{Ԃ�SHk����6:G:8�Tc{�\�r8GM5�5u�vē~+W�՜{k����:r(���)��ʾ����V����z�̖I��,'^�*
��W��I
�3�:nJ{V����;�7�X�1�P��S+ny�>���ł�T�'�A.w��O>u#_튃js$S��=țm�hǸ�H�ї,i���8P.���u��z��;Ǖ��1���y����R
�4�����c�ժ!�
m�����)�վ�:�Mf ;�$-��]ǁZ��+1�I���������@�4�G_��EQZ�J%��9]4)�gno��Wŭ��?���<`�_n���6$�hg\��ʁ�|g+�7�#A���{z� ��`�D1�������%Ȉ���o�:�t�Ȳ����&�`�{p��tp��Z�nW=e�ڥ�N�����K�L�8K�أu�)�9;O�R5�Wp`�Q�Ǭ�r����;��Sn\N\W���h<5�R:�){"�R�s�6�9wC��h71��/�ĕ��v��o@y�#f�Me���cV�g�4�Hp�<%⨫�m��q��8/`hɥ�Hb#
�J+hO����nxP淇��3r+��p�,�����S6���N8~��<?��
jr��w��s�bL��r���^J�
�7�E�p��1�E}����BQ�F��춏]:d�zQ����xZl�ю
���&bbwN���w=�r�����3�Y)�i�>�A�h�Y�Y��+<�Au �O��}�j/��ė`�#%��W[��������.Ҍ�~��F�a�(^����ʝ2�>��}3�:k�<u�Hp�ї���A��y)�GW��{vbq-Irt��|�츊���^����v�=ٸݑ~O!��1L~%��&��hjR���
袭�+9C���'�����N��a2���W��G�i�0T�߇�C�EI,�釼WN�(��cP�7����&<ad�n�w�En�<|�e�D]�'5o���L^��������Si���C��a�"x���ݻ��N����8j����K��\�QrѨx��ڠh����8���I�G<��B�^pҜS7+L מеwV�~��V��&f�F6�z�(��1��T ����d>=[=~��!;��b��4��n����0�#P�/�����ƌ�e���nF����E� ��y$!��|����Q�JjY������I�(ΆƏY[}���.a ��ϭ�bO�˂��\�h��j��E|=Lح�P��3�����ڽrUsO��R���ڑ�rwl��!<�V��ϝ�G�p���� �
��N1=�y�����Ua�����)5���2� �V�0;V,v�R9(�����Uݯ���U�|��Gw�yc�V�#S��x��)�K��w��{�.���i6`k��(�o	]���a *(�O'�8c�x��0�g��7�Dk0yf�`�t!��%d����i�i�����Q❧�c��҄?�5q�D�4W��3bkÃ�� I�/�P�5�8���V�G\�&��0��[�5X&ۧg�i�`5xa3y����5�R:r�oք�e�M�E����0Y�!����XX�"�S�qaJ�z]<���b��šJ�@��MS*J"йk��#^�OtT縲�� ��>��H��+`���A��L�߱p�:yɸ{�| 6S�#���O�S���-�s�h:�S~����J��ɔ� ,�p#|���XX��z��],q���������C2�h�H�ͻ�#��Ͷ��[�O��K�,���ު�����*7F����[���[��8�V��������6��}��a<L��Ԣ�)�5��<b�'"�hJ��d�ot�}�����J$B�X�@|�K�N7����8[�p����E�Y#���7o���=�(3(q���\Cv���?,�<�������SIܘ.������0�#�N=�!��|�_��t[�oy�Z�)���T��9�H]cu�!M�ce��Z0��stLx(��#.��*lMH��/Z�~�%��s�-��fZ�%�}D�����T�֋|B:�,�a�"��"�Kbo�\�)�?���'�A��d��ƙO췐�;?�N�3lA�\��؜5��t���뚩w��m<���t?�N"�/��E:S��	��yKGp!/r	U~C8��χz�$5��HQ��:L8�q�"��n�;i����nj*27à�e;���Tn�?��j�@���>E�++]I��ra%���Y�X�x�`Y�|��Η6蕣-]8�
�}�#h?�YO$Cl4-e�1��T9l�e��5�������`��[�u��6>�@���hi�w����|S@\�̙S��)�W�4JØ�͟D2??߱�au$z"��D楎����Yo�}c=p|�0{�ȑ/�>��{b���Y�U ��i���Wuk��4�{���M<*ep|�s�X	3�u����e��{@2�чr�4']���SxcK5�J{0��<��oL�����et�ZhDG�%�M���!��� �};��B��8�$j������=��,~Z	/��g�-ާ*��Ӊ�ȘsP�0G��!�J�K�hX���`"�<E=�Q'.N^h����°|ˉ69Z�(|(�ٝ��M���nVU�� f��=��q�ce���i�E���KG�c��m��)�N����F��b�Ðۻ��P�Y.�G�;���2�T褀�ƩDG
�1��$��-Nx��+CtR#?H'6��F
g��,Ԥ�1�sѽ�}����0c�o��4�4��Όw����ֿs2V�G�	N��5l���l<A����^�1/�`��z@c�qPe��W�8$u�s�뤩����VJ1��1Opi�U
�T��Qh���w���v���5{�#�^���B�!:���$9�r�6jl��(�BG�J-���^��%Q��Sw�ɵj���X��	���q��ډ��e�f|�HUe�����mM�Z�/���u��+I���i�վ����M��	No��H{��(�/\+Y�/y�W�:4��g {U[蛔=NtvIU�"�N��$��|��(Lm�q���T3��l�8��"7)���#)�m���l��LF�5w�B����NXj��/
ɷ�r��D��CY7��\w��f��-(���nh��Y`��t?
�b��OEz����M����|�l�X����7����h҉�m,o��o���9(0��f��j�gL�@B��.+a��Q�sOe�q���/ik��ᫎ�L��{�Z����g3RA�Oy�0�e�*B\.MIz�bfۦ�@�����:����6���E�L� 3rm>�{�!�Z�0�9��"X ��tk4Q Ԫ=�U�_E=cW0�Q!��0b ����Ȇ����Kb1��p��åN|���'��hy�U|��/�ᑿ��;!5���C�z�M֙z�:C��T��_Q�:���)��-
�d�pN�F6O	�t�r����,-`�ʬ:Ȳ��:�	G�ϖ*�f�⮫W����a�/���)��v�H�G����P)�Js��uAZ��C��3aٔ��dr�^�O9�S�UB3��	yk�&Bnג�����#�$jT<R�ʮ�	E	�d����JO��X�=S3l<.��6?\%5*���"y��dq�ۈi����y7GI��,$ �(Skph��-6�
���`��bPZ��h��q�)LQ��`�g^B�-�2M���I^���; @��Q��:ވ�C��Xj}s���|d4`J縌����fY�ίaXֱ��"�B�U�}�ġ���(J�D��9�7��BM>0���������u@m�]P���Th}��Ai��?��[e�귕��� lE�D��j�,�FW�-��UzD�fy�9H�NOc�hL��FG*�f9t9(��h���)V߼5��Gˮ�]h�n57���_I9��y�9pv�1|��U5v�+S�Є����#6D�D��%���)b�ۄO�Ùտ.��	M{�s1�/��6�%G��L�k�a�F��9iC
6A;([��u�9-��0��5��gE|��=YE��筺�-A��m��⤶��jt�j�/�����ce�,�}q{�]�.o��&�W�G���\S9�`�)JԳ6�E@��^s�a��<Ѧ�P��QԤ]�7���<oJIX�T-ַz��혷<`��-;��O�6c�=)�ފ;��n%2`Q������hP(z:x�k5���ד�_=AV�_P�z�C�؈���Օ�p\�i�mˠ�t<�ߛSP'|�{��}��*�&���UA�]�}�]@_Y1}:H>�E~R������s~�gM����{�+̉��ҿA��}�O!�\���y��H&﹅P����V�C覆��I����ғ-]�/S��˔���䦴a�oBC���42�A\��]���t�8,��[_�����?$���b�қ���^�׫��ߵ/���. JPw�,��R7em��'9�_b��`@^�Ru�|o�Uj�|q���A ^�.>sP�v��q��4n�nH�!�=��#�艖���?f[<��:�*W/s�?�m��!׻;�
Z���@(��妽�l�I��
ƚ�l��{���z|^db%����+��p�� ��jQ�u]��F�D�B�7�<;�n饤��r��~;��i����ay!���6����d`ډ�+��<υ���ul��&��# L�%�[���bt�\�]:�-1k��/��IDX����xB=�^��0?�S�d7�Ν����C��b�E�>�}��0�;^���`^O�.�B�N*�M#WB�G�[j�tX��6���+:B~DW�I	U�n_tIJ�R3��ZogQ�ms���J�������1�f�L��Aj7v��\a��rz���q��2x�)#�a�5��J;i�mB��"�]�t�n�{��מq�qà��q��\�_�����mn�7'1�N�z���M:��=g ��Rr��.���S���(R��],8�&]T��1ƍ�u{�lZ�P��~ M=J�/��ľ6'յ
w\z�}���6�������~1�I�&X�"t��3��e����J���ַ}���J!��l��LdGܷ4�N�>�x=�D��I�n�/�c��M�j�2V��*?��Q�Lp�ؙ�A]�<�y!�����[�3W��]J�� �������Zv���)�]Js�C-�V-��0��Z����{\��ג�t��U`;t��D�n��C�l�ؗ81y��X�/�������'ݓ�<�Dm%��-t�8��D�R��S+��iF⌗>�YWE�	W7�7i��n�K��!
k�o5�s�)��40薷&WG�-�2r~�2�� <\��I_K$�T��و�/��B-���i:�i�ò)
r.����<�D1��	I�LQ��:���}ytR��B�aFb$�T�k�A=C/����)���vl�ܢ;�G!�)����2O�S��Ll!J�2|.uH=�ŷ7�DE;4;9�������;����㻞ڽZ��<�ή�ù��[�,h9}>�P	�G@�H	J� ��M>�n������I)�r���_-�W!��l�:#�Q[Q�|ߘ�ҍd�_�x�k-C�
�a�`ۏʧr��&[���&�b�_�RZK��"MX����G����xO�ݛ�u-k�=��]%B#}��~v�o�I-��r5M�JZaï�e"G���v��ś5��;E2���<�, Q'�bл��:ރ�j�xe��DV`�~�5C�'�%Ǩ��ϧf��[��dE;���CXC���~�{�s�1�_����N���8	��M��˷�K:��#z�$�!��l=��%*���7�&bC��HHm�R�m;olgҸݠZaE`nTq�MQ���9mT88��v#0�f�p���\��(�!����*���%�@�%�ߑf�ե4R҆9ޟ	�����X��C'��8�Tho�_���-�J	�e\b���؆����XK�u�7ԃ�2��5y��같��<��98Ză����"ȡ'l�[�WT\�u�%7�};f78�'���H��Ū�( D+����F�W�):������*�9v�H&I}r,g���[b5��#�;��0��f�r:Y���59,�:v�p@�����s��X�^N��d���u�j����WH7vhSm JJ|Xƍ&,%,���z����L�=SA��1�Β�Q�۽�zw�B������bj�b{�٧ �{i�؅��T�=���PFC��~����W��2�4?5v>��1��훛M����o9��.�1���s��>}��~�l�W$O`Wb�W��p*�q>�t��(JWXC�̠�W;o�b�O�nٽ�]�^4*�x�j$h�}�3k���z4�,e6Ė#�����A~N�7������yVS�=v�6��C7���p�/�?C��U������h�X�g���1'�1`�pT��V���.R���|ŋ��ϕB��$����ފP�O���;����~�ww���&k��S�E�E#u�����	�е��73��L�'6;�����+�+��j[���t0�G�??���u��8{?/��������ψ�0O޶�Li��yL�q�M87t,�c:�Cn/�|+�}��K�S4�x"-�Wk�,�1iKŊ}L;�"c,�R\���<��ְ6�+2����>�tX!ƦL�}e�Ăn�d���:;�Z���a� �X����C�������?]m��^�
�n����b0߯��[r؁��� b��{��� Q�ɲ����e�P��⥳w�{v�����1��'��>�V�jvb�樂��/oBC2����d5°A���L����hhb瓉2��g�)�Mω6�-KH)~b_`4n�k��5~�����5��UO����\g˴=k
��H]eBxۮe�/��%��H���@��rV��jW�X@�D�.��ތ��I��8�������.�9U{��M�L��F*��9���i��Ч�U�N\E
A�|�nf�S�+�$4����G+o#��z�¯���۝ԋgȫ�6��%:`)\|W�NŖ��Se*Xߐ��!�0G��'�/[�Kr�TSA�mq��/�e��f�@�\�p`S���ؖq���G��4����}��mo�����:�v��Zw�-Y�?��m!���}�.#*���4�(�)���P&�`�d�S̫���C����U�V����fa`��Tz�����W��=�eNt+�o4�V"(z;裕��)!�mF�������bL/h���Y��,8!�.�ήV��0�V���w����:���* ���*�F�|�S�hIG��Ćd��c�I�T��/1�ER��+u��\$�iV:D�R��A&zA��o�8�2��������e30v��;��T�)�8��7=�k�B�X�4��ڨ��9��Y�퓎���P��&$��`�XX�M��?��}���邤���r����� �RWD�Q�x��âZW�WM�ׇ�)�}��`�l_��������ܟ�Pm�\m	4���9�z�qe"=+�6���7��f�8�셊~Fjr�cJ%(sh��W3{\N��1�)��O�VB#��JlT`7"��A��u�;K[�,uXD���zj���7�3�0(�
@SЀ��r����dI��yG����L����0���س�8[�aV�~,�j@�rS�W>���۳J�(q�ޙ}ş�b�6�R8qG��?��x*�c��Y����Y�-�к]������n�rۀ�pq�5��<�~X8��T���4ߤtU��0N�`.�LI�~�e0X�8�'�:oAm��Ǘ���
�h	���3d������2r�6�M�]��$��#i��3nz)�$�j3��*�T��ȭ��(��,������;W��Z���JI�5{��(4�2��	i7�	>Cb�l��4l�$&�W|a��o�}	3Fjt���b~� ze�ι�=��J��2ƘX$�4�,c�Ll̳��e�pp���������5�Е鍚�+�N�8��y�7/571����"2�*^Vk�umO�p�>���`I68&��!��	k�X$j�y
��xk�V�xɰ@Nrx�U9=ޖ@�4VI�����9Ҧ�`����0L����K��	�둭�h	["hS�&A��� �޸G����u���{P���T8��CP�œø�E�ǾV��.0e9�;+�ٕ��W7٫S�C| �V5/\�n��--z��@<�Zɥ� �U���Ab`�̣�H&��Z�Q!iߢ�U
�.�A�l�v i�ʱ(�
�Ǭ�Ν^}��3���N�>�<���t�74�V-��(���$�y��2�=`�kv�*��<ʤs6�����o�|� ����c����g�D��a��OAY͙���:B{R����F�Fܣ�DGAMSI���@�<���C4EsU������b }�7��M�jp<���xV�PS�������%��>&��7�.%k��J�y��48��W�`xyQ�ᶉ�)�1{�>��j��XӋ��T*��h���;�ө+JCQ.0�u�)`%��2	#�a����h��
@Bz)�d�ɗ0�`t�R=m���|L޺�������Һg�qY��u&�`�`,yτr��s�q3�}��(+��y��P5������bT��j��}�;�67�`�@�,�<����V�ChPtÝ���Zղ�1��e� �%U�K�(������N��  � ��@(X���qRהQ�xb��ِLB?S�'�*������q�$AS�f-�����B�Y�.7���m������������ ��XN�"��z�O���w	b��� �׈.g��3��K�{5��Y�%[�;r�'� ��<�A#ñvj�e�,.������<Z�y�xAT���䬤�P_�=]tm�՛� �}[J?����Ri6�*���IΩ=mC� ��F�#X��*��p:�^�T���[��_���Mg��`��#6��)��a�N�ƛ��P�H'~�Z ��c�%?���Jc��'�Kg��k@A��Y��%
�2:׆��Ɣ�����H�_�FoQ�8��t�a�6E$@������,aN~����Dd);�k :�����d8�9i�!`o&:���[�RK��[e�1�;�13iO{���"lOB���U��~����L���^�����G�m`>=l���4!���-�Yk`z���=����(!�b��cn&"��W�*���(��_e�Yi�,��_2�z��޺r���0J<+�oD���F0��4	� ���g�.�^b������ipД����%,AQ����M��9�1���^����F�Z��7�j0*|Ino�U.��mD3c+*0�E�Jz�zgr	+��a�^MȦ����4x��*.�P?�ܨO����E��K$p������ћ���K
�k��*�����Y�,�~��/a�ә��BS���rd�m�GPȼ�����Jz��]�=�Q�ߛ/��hL� Ɵ#n����M�X�� Q�w$ �<�~S��'��1�v��?������<7�L"���ZDp
��v�/}LX�� "��r܃��q�rE�F~;]��;�فq��Ｚ���ϳ���k�@5��K٬)����6.�;H�G�`��"}t�W�:Wq����v6-�ᴋ`�����$U�t���VQ_P:6���7�ǡ}�Œg'w�Q.�k����~ݿ'�Dm�2��%ohU)��T�(O\��������55`Z��N�1�wPVD�H�^/��۠�n9��K^�vM�	��B�g(�J�A,깕<�7�F��ΪJ��Va^zR����{���H�R�?���k�z��V|�u>�5%�o<H9[�LU�Y��NF�����R�P�q�Z���Y�'�l���`��>�3H��lh��v���S!�r7����#Tsp�BJ���!6�׿T�{�4��������p��<J�'4�����W��+��ʲ�+�����[�JA�(�'_�	]���fy,|>	*l��ͮ�[s�����K}D� P�%l8#</��߁��up'��(�۝��� ����9u{�Z ?��zn=E�m�\�I�up�z�m!��;���\�0y��z%-��tr;g��x'W�޶$T͙+�HD2�	J��4��W��؈��f�L:�5�\䙮����$����~�h ����ɝ	8��ws)��)(�vBHĿ�;X�kښ����(ck�m����Z��"Jb�!�|��A������Gſ��j}��(j>V���-��P�Q���7�˪�nޏ+n1l�.��cQ��l{iZIg���7;��||~Ƌ���4��C
��
}�m���!���H��N�H:��)��V��֒;�c�Y�B�A�Li���[����!�ֽzr=ޡ/0*w���#�W�wLw�i��\�����rJT�O�j� �W����'e؈y]wx'S<4��։��i���e��Q RW�{H7�J+�����ބ��+�'���n��®u-�-�f�Lw`�S��z�����(�O��\m�8�N��32|��{�&ތG��T��� �q�͊�S�����4��R�)yq.K񆺲��^��B�*Z� )k�Laf�$�\?�XX
��3��E��A�����Hj��[ՋH��1iȶ�v�� �ͤ�T�=�����y؊�-��V��b����ya9�@K�Z�|[OT M�BǾ�D��z�csX�_����O
���S_AL~�D��w�gi�q��/���|�7�hc������X>~�u�x_ݐ�M��ۖ�C	�n��{�h�Z��1ᩎ��|DS����C�_F�o)���SmÞL8������!z��iT�Xճ�{ss��W��I�>��.�q+����]e��큏���{�b���R!;L����b�г�����.e�L����!<�����$^*g��<�V�yq����x�3h���VsV��#��	�W���g�|�IR�!�ļ潧f��[�ʤZ��NF�*Hu�F�%5���([#��r\[��C�S;�"4L"U٫�,�C�T`O9���}(B�:��Za�A!��G>0!��WD6^n�rlR��R�K��IE�J2Z�.�4��J4��\^U�4;C�@%��(b7�.^���\���> ����9��o��;/�8�0�E�
�U0`��#g=��
pR��gh����o#�,"��6 ݽb�3TJA��rr�o�)1ܼ��9�O�d+�YL}�33�D��1�V1Zߦ����W�� ġ�����~��r�ѷ�*f6y�"�u� YJ'�x0�x��LMVo
�� �EGTwKx.J���%n
g��v��%�|�Γ�=ʎ�_�:���K5�m�&��/�z�b;�Ϳ����]qye.z������n�m#�B���!T<�Ez:���DI���/��hMN�9"ȶȖoB49N�h_�o�:%<B��n3.���QCqq�6O|U�=�X�^@~?����\���.�(p��'�K����]8��TJ(_?�w�G�������	_�Z�̋QqYH���ဨ�!�W��"ݳ33^K�.4e�����\��Ց�f�>Z�
Й�i_B�H�U���m�����Z�Ɛ�?	K�&o�@;4���e6Z�8\i\ɻ�R��3�����վ;�|�V�!%�)�*����J�Jf��A�8\�N��k��BׄX�Q^s������@�h�]�64���1�$z&	M����l��k���M��'x�j'��{;�tf�&*9-��\&�:Q��bё��o��BŞ�9
1O�P���~�H��sq���
�����1��>M�	�܄BPȞ^`�\֪h�)K'O}|ͳ�Y6�<���#is�Z�ɰ�8�ӞE 5x�p��q_���B"c�5�{�Nw��/�����6D���_]�s ;���K}>�i��#R]�~��n�1H�e� �1/|���#��2�-7��	�h�qEPn�oa�.�F��Ϯ�؛]�$�i��eO�?H%�M��ˮ�J�N�`�i[t��M��jA��$$+tْ�*`��Nb�L�m�li��X��N��"�����2�5���0(AN�k�BH� L�}�0��-�??�2�����5����ol�������g`���I8&j�h����:���w����콙���b��}�U2Q�lj0�yX5���>�k�2����u�*�Gl�-�p�iq٨�lԩ�z��#����=.{�?��- <��x���褚�4���N�hc�<2-it�xCI`5�Ζ
��߮ ~ђ�܆��e2�F��Ċ/�6ԙS^���t�[CU����-QKW)�4������mFŮ:�<e,��ka2RO���}�/���2qGRIP|t08�F�`�'�F+�HD������3�ԹP ��q.h��dmT?�#^`���~W�Ĥ����:��nu�zִ����&��U*DN`\�&W�w&�5Ԣ6xl��~���4Ƥ�MӉ�c ,7�E�����3�f�I[�r\5=���
'`�@�/H�������_��MU�TR2��U�4����#�ō�&7W�m�Y�IK�[�����I��j$d(���%�~���i&�M�$���;����������$�4GFZ�0HY��Z*DD��т>��h�����)��ꔪ�='
$4�FQ�2��"�4O�x-��<N�Ғ���w���}��Ŝp�;!3U����������o�s�0��U6a?%^���*r"��b���i�#V���C��׬�gn7Ie(�2�n�w���|`m,�哲���wL^�pr<�sb|"��U�-�mYW�|���۫Q��m?��F�JtL���~�|�j��U�e�I�vX�nF-�(uFk�ꯩ���������)�J&?\G!功�D�S�9�r�o��)@�0L��2;�α\���E�}]�hQJ�޷'��p~M�q�C2CΦ�#��;m ���˟��2w;��(`���͘�F=��'��Դ <��K3�����yu��#.6����+�P�H趱2�q�&�y���"�D�|�b2���`����*W�C-�B�tŜ��)�� a��ԯ���[�x�����i#�(ZT�b)"q 6���-7^~��k#����TY�(�fχ5���O.�AÑ=ٜ��o�[�� 5n�/�+�EU����b$Ԝ�n�p�:�LeU�&�f )ڬ7�����4��r�H�Nt+�xa�G��kb50��@ߞZ)�y���Oz�oTX���+Pm��t�@�~���,+���Ϟ�Yb���I0 �sU�D�E�G�I*&��V�ڻi�ѧ���_dw3f��8[�<��7<w����aM�*��J�X�?��rr8�V1;��;9��%~?�SF��OL����B��.W��.мh���κs�֞�247�L�:�m�qv?�	P��6���ZZrD;�;�U}�]�~�`�����P��EUy|���;Ni8����I@�~?�@��3~L툊O0�0&� ��h�b��k���q��4�,��U~W������r h:�\w��rCڧ�X�:v��}�����*�ϖm�JF�z�	E����Ԗ�9oUj:�|���o5» ���MI�&'G&q�6�KC����}��Zո������2����������ݜ�DO���������H6�[��?j��Tu󀶲�"o@�B��M�i�����A{���Ȗ%�;[y��|��۟��M�u}��==����5��;�wU��Ϡu��@o�Cv�"Wr⭰OV��_�b2�ӯ5QT����oP��5�Ə��;�8~Ԟ�[*¹����j,.�@.�$�0�S1����S��f��8
A�:�r��AVq�@ɞ���	-�I�, $AB�?��^b�Z� �V���EUc{/��e�Ek��]?Q����V�!#����±w��Y�Ü�}�uˍ��y����lA��Lݎ�ח$j��`&�N���@�%�'a�� m�����۬ϫ�|�ub�����[D�8���i�Sٽ*����82M[+���aHv���4^5���I��G���ļ��j/Z�A{���\�Kq�E�7�\K''MZb���:&��Ζ����I�������Ķy�Og��-h^+�%�<�������7n
ku?�i@$j��?��J����J�t�+���;m���V�j� ��P4;������oQ� Q;Go4(7�'�&_Н吧�������D�-�����@-48�m�>s�V�?9����Թ��
h?�`.���x�w���v-�#u���%���ֽ}�Ju�����h����3G���� ��c��؃~�o#Q~%K>�n�0>�����v��$�=��۹�Y���s�o�-~�DLԳo��j(����J�f��0�ihrS�I�f��	��D5��e)5s��O���H;��x� ����n���&��҉�j���5���3�8C�-�����N댳��\G��޵@6P~�:���9��'�mlʯ�$��^��.q����K�����x�F���.>3yu2,�V+���v�Y:!1�VP3��L��xY�M�a�F��YO�,y��g�F���᭺s�3��M�-��yw�8{��w|?qJ�4�HO�������q�c��k�ToP��f��eъ�ϙ�ANjz/F�����m�Q���_��lj���?�i�4�k�i"3�U-'�����u�؉�^�/�j_IʧJڪͪv�,;��^8_�f6j	����t<M��������H3l,�r��Чr�(iE�ƪh6pB�Q{ր��'������k ��|����8!=�+�=�?��F���(���qq��x��)Q�x
ʂ�H]�mlP���א����Mq��<#��7�{>�ć9On�����p���$�zBC�>�Fu�Mlq|w�Q����U�։�Ts���C�Z5��x�Q_?N��7���ϝ?y�@���[�2���B�u=J?J=��k)�O
�$��:�-���?0�*����q��w�揕`�p��(��!h���T��h����UiYL'�����P8�����\k��P����ᆫ��?�	�d�p�9���*�R
Qa��Y����ȋl��\_sDSÛ�q9>�T]h_,]��Dq�F��1Y�-:�v��6e(�S����E7V��u��3��x�g_{SN���b��4q��	�0�ك&j�-�^ʌ��m;��YJ�a4:�����,���I���'���>��v�������3�=;to�z�z�������P� [���Q�s����.y�$�?�;Bab��$[Av�.V���,�Zxx�����w�<��7�B��DC�O!~�B����
5+�l���`TuS��[(7��g�m�?��o'bl��1�vZ��XX�l*��J7`C�ɾR��â�s'��B�1�E�~�|�c)��e�g%�H������Q�>�1�y�¤��hoV��wvI56�@���z�9�)�"?��1ʞ8(8l����J��Jy_�7�o&��Z����j��B�?����)��0<����z���Zv�x�-��AIW�Bcw�#��&S�]?�n#g����{�5qOm�$muҿAW��!ђӁyJ���ɆTt𷈑�A�#*!"~�g�u��<��n$S��Xd�1�I�KFMҊ��.��yN%��p�+���"�u)��5#��t:w�6�.��ƭ��i�ɩȘb��I+{� ,Gc�WD�5PT���_�n��J�	���n w�CA��x��mGrfi������f�U��EB�)~����:�$%`2P�^{ՙ4^�� %���5���	��3����p,���%�rP�s3�'V.�󢇁Jfv�3���R�&�N�����H�'��$%L}}!��ja.Nj�wƌEJ*g�!$J�jO��ܒi��ܿ��p�y�rX�)�R�"�C#�kq��8�\ ).�c�<B�Ӑj4ԎV˜�N)!Nx�x.���}�g���C(�#W�â:����޷�����O�HC_w�4�$1�����r�N�C� ��U�y���A LR,�$�Z���3V���C�Uً�dͮ/D���K2M��O ��t�b8峹K��I�f_�9��X�7$ٌ?�m�FR%/L�}�ظڊ���E���Y����)�<�&I�b�����*V�D]��3Ğ�y��U('�v=Έ���L��/H�m�>'+������c�S�R��M¢��<2�e�n�����)N#���^_Xń0���-�Cm���Q�������uD�W����gy^CK���9�d���a�H���P�̲��Ҳ=�Ά�W�K�Rd@��m��	��_��sZ�X@�Mbtf�*��y�ʹo���.������Lշq���(b��^m��>}˯r�h��{����!��i:�f{���"}a��}�S�|���N�9�JzP��[Ş��q(7�t+)3�n=b������.-�E6
��UGg��;ۻ�VV���l�m�� Z�-��%�J*O��o�ٚW.���W�,V�\A^�Q����2��C��5��EX&�"w�9��m��1݈E��tj�OZe��&S�M_5��BF� �0f�M�5&�xb�F�.`)�&�A��
��]�Jϒ����{�� \�6��CD(E!��d7�W�su�K�s���:���aZ�e��CΙ&c�(̚k1�( ;�Z�8j�1I�6�qd�k·���5�!G��&095�[н��`�^����
D��fF��:K����dc�]HJW�=���(Qx�{� ���|�-��>��RWX�ݝ-����u���$v���Ď���%���)�[6��~��y�J�2�6��d>��)EQf��ϫ�ƾ�?�k�[K� R�>s�bӷ��J�ƒ���M�^uB��L{�7l"�~ǫ����8�
�qĩ#X���G�B��R��H��a&��)/c��~�I�&��k-]1/;�R>a�������{zT�k���^+�tg�̜E�T�מ!E>���0,�i��ڠ��Du�0�x�YndxF�x�~��qz���dS��ira�*���LB�/jw��.�g$��F`�������G~�R�2���p�����/m�7G��O���j(���p3��m*��~1�4B'���H��G�_��̧�e�w�c8�l��rCz�1�Bf�2�H>g�E�]K�a��oU��,���-:hT��a���.���H^zp�X`,#��r��\��=K�J�w���Z����̽I�,�ujQv�q���5)���3��+�]�G�qT+���12̉$��9d\������|ю��^.��Q��P��$�Ӵv�eq��l��Bގ�1�\ZYXH�:��8�&H�s���_~���v�`!���hGD�>��C�`fN�7yD	�tpO��j��4r��_ܟɃ�ؔ�z��+�\�DՎ-v�(5��%C�5Fݴ��!_�^��2�d>�>�x6����������� ���	�b�X�؛�q�����vL����*�;.��sd�[�b�+3X�#�gM��!��%���4��b���>p%�t>�-��������D�Sl��I8�j�x<~@�zr*Ky�gc~�����c� ��rԓ����v-йڶW�B~����;[��y$�H�%ND	~��i^Cƍ�G���O-��;%~ZP8K�������9���F��-���1��+^�jӟ�U���S ���u=�����)��8����+�;ۍ��bDs@_�@f�`Ule�@���6n�7'P�\n°r�uy��D�O�S�8�c>�q�dj��6��3VS��\pֺ�Y��,����^kv��5wrH �`����+,#d��FN�4��$"�Įt8)@]5p:H�jv��R>.ԅ\�:?c�����2��b���#N�Y�����5~�ʄb^�$�a�9]~U�qX0Z�l@^^\�.��F;��7���_l�a�xcWW����.�sNy>@��e���0�#tO�V!��?&�b �O��i�%� L$�mD6yn�����\���M|�~�72a�9�p�G��`��x5P��O2���E��WQ�VQ)��<���-#������R[�__���L�)˔�ɍ}����er�i��^�5��ܳ�ʢ���)��/�Zaп(�ӌ��ǒ�
q���@�Ǻs�.9a��u<F��D��~J�<�{� 1����y�����nM��d�&��<��[h��۰��,�� �#�F���WND����K�~��� ������	!�^C�*���LCO a7��#��fj������[~���G:ֽ��~IՐ�Ӆ*�
A�Z�}��-]�����ެa��f���>uQRף��_ѵ@r��λ;���3ѷi6��-��u��n���T(V�d��k�;����ӂ���P/u1�������v:�q���ރ~kj:t���l�O��?��o���.�Sb�$�`�2�,V���]Bh�}$A�\%�q߻�A�l���EU�?��: X�Z��.�G �}J�7o��8[��b�(.H�:U#����d��N#�Sg��w�X�}��٢��{���d���%(��6Y-!����(zŅ�L{�Y�d�L�:2��'��'��`�[��c�ˌvZp��<��3�;.5Y�G߅=Y�M+عU����+-n��8�����`V3�e���:��(Ne:���S��!��G�>դ�c��Y�E!�5H[��F�T����wPN
���^K7<W������1�?��;��'e��Hz��1�G�յĬ:յ��g�PQN�4��E�!ѡ���`2��cB�� �!��O�`����u�Ì^�I���1��##�.�!OȨb)YwҠk��d�c����LGX��U,â���`�`��|�BД�W�C��w:'.dڔ��-AL��	�P��d�lV�N�0��(Ջ�2F8�d^��FnO�T ego(���h��H���*U0�H�@,����7�/��#y�eS��K�76BL��͠&��0�^����x�L�A'���%��h����z��X(<=��/���r�'���bn9X�C;�C�_��'����-��ET
�xԲ���h$[ּ�jƢ��l�������ۍ���(���8�o��i7�!v�p�d��>�+��-|i_�xd(�����Ù��𵽥�9��~� -��tu� �zo�W�8�V�^�n~��k:�I+Զ��X}�ihGE��u�O�V������)�{�
ޯ6S�K�BP�'�a]l���d�װ��hҝ�*�&X�%|�f����ՄJ:�Ӟ�JɥO�"�.!o?P]ݛW�z;ӧl_��F��0}�g���?��,�45����+�?�A�'�0tF�h@p�쿫�Գ�df�����B�ڸ-$>����N�ͧ�z"�ʶ~��?�{��8:{���c�׌D�V�LP��d@{�O���T�ɩ0x��;���"��c��}��*��e8;j�Z��9��qk�-���N=Lx=T�����_~��oS_��a�~C�d_�g
�k�_���3�w"ud9�8���{�E6��o�V���֛M�R\���T:����!�j��B�h�	W۔+�m�=o�������p�b�2��a)O�v*`��X�S8ٳ��irO��Qď����=���8f3'困�b�,k�Y�o��X��z\�.�7�Gа����)\���ʟ�v^4��̸��ʋC���3[�4�!�)w��J^���_3�	t�xɣ��X �����;�6�S����::�'�c��B�B�:+ʔ��r�<:��� �0��$U�Ϝ��0]��7�1��`�$ڌ���V���.0�%G�Uû"�t#�#�᣿�.zI��g��Q���O�C���&�\dЅ�����ԡ�7m@������&�KG���M"���tK�z�'R�l�?���4F'}I��_�C:�����B ]��'���z^�A(��?�ʋ����A��,�Z����iBÉ4��@ۿ1׆Q�B��aѫ��;֩}��gމ�~�R04��}tE��1�����Լ8�o��^h�s�h��W�@�s�����7 �E��S�2���n�}�~NĲ���j���2 B�R�m��4���O36����y=���2��\�'��+�����ҷc(U��g�ҍ_W�j��Fk	b���W�H<ń�$4V&��n���Ow���=|6�l�_�Pαd(�l`��W�E�5��;~�HɈ�0�n�|�QU�ݷ�6���0D�a��M� �H��.�"�2�b�rr����Y�E�/ŕO/�E(]���l%�hn[5��EW
e����r#��v=�j��+8ʚ�UFҾl/�P�.�G��h+T0!�J�l1��~��ࣴC�U��e�7Ht�R��U5�����!:��O�S��U����j�i���n�љ�ń��.�7�@u�H���K�}�Bj'��,��[y��kȋ��Dʭ_4#`��S~��'B֋rB�V΄%(�c�4�F>���D�֡���z0��Ț�g� �c�x9�m��%�_�-Tɓ�٬ɍ6�)U���9��T�x�_sq��˃�0R�=q�KLK�&=��aP�|$2���ȩ�_I��%��x��W�4�4g�yޖ<~����l�@%��wh�v�t;���2�籓U^df�pB%|r�{�t&r��c��u)�B��q��`D~�'�/.�d����s��rO+�y�j�}s��deL�������b��3�ҎS�R�W��['J�� �P�u G��w)Hv��P��u��ї�08'0�� `�6;��{L$'�E|� �=P�'@)�4�*�ȱ��9�ݿ�"Z�]�U�A�
�@@gl Yc�W (�^k�6�VwA^��]I��B�;>R��N���6��fy~Ѱn�-x�u/��xk���7�Mʢ5��j����d��i�8�;��n�-��
ck�:��9"�ܭ�d;� Ӯh�/1"�k�F�s�7���՛q��]����#	���iq'3?�5�Z��.�u��}�߻�K*ٟE1�L�c��@D�d��l��:��:_�s��-S�5��އگ���_.��?���$��[I6�3�����G��}��&��tҘ�R0�m ����wJ�������e�k-��߻�9�o��aF,a�����s��
���NO���t��RN�u���
����r�0ԫɣf��}a;r��l �P��q�i%UB O�(5/�x�
��3��͞������'�����3j7��u( {�g�ŉ���ZG��|�"�Z�sH��#F,��NP�����ᅶ���x˒��2;>�K~����M[{�m��7<:�o8O��3<��y.&w����X���V����b��O�2>�p��۬B� ���/��G�6�.&sd��,�WF&w�iR��c��a(*\2��@�P�̪G`��o������l��`D�S���k��X>�R��z��i��u"|uz(U<��#�S�0�|��YY>y��'�3lI
JI�U,5��8#{N!Ж��~M�~�������\���i�_�U��o3�G3���4��by&�$cZ�r��QI��T푾<sM�&\���A�ٽ�HwU�0�~f>�A�w��@&���`hKʾ�܏`��=Y(�*�ա�Yſ�o�\��s`�NYұu�����76;;�~�mE��+�d�-�L+h�uȸՖ���s��`7�>��]?�{�L�������;�o���A�xm����Ü8b�QqxR��\u��>(����R�I�G~�xh��j<�^�+�2h�g�ֆ�-��3@B-��h�䁹'(g�JF~��fG� �.@�to_�<b�E�g� ,~�H(u���� �Q����l����K�����b ����=����Y��X�s�ȱFf�d���x�i���Y�D����� J�\I-4R�������J�^�h3�������,8��
-��Ʊ;��:��j���M�\էh����x�ܻМ�y�:�4�zD�.Q�sP�KOr��+�b�Y�O��;��R������������w�TMZ�(�k7��=��kܟ�$R����և�͓0W�v<�1�3"I��S�c!s_ih1��5��H���վ�����+"m�$fl_�1lE�-�u[ �^u�~��L� D�V�Z��vR��e�[S���a���q1�q���v���E�8G�	m =uj'�t��m$uE+M;1�%���}���i����e��Ņ���#5o�38�E~�K��uރ2=�2Pck=����d�������ʐ$�����l-'k�_d_�֜q>�'y`��2&ֈ��=�=hk����T�&p�����b��.F԰a+D`�Z�P�Ӂ��4���R=<�g�x��eA��g>�# ���Y�?K 6�_p����F�|�j�	��N��R��cɟӉv����:�� j�ğ���ĳs�U��Vd;��Ɔ����G��lq+Tn���h�U���"������G�P��&ǐk��.�yLҷ�5]��-�[��Z}vz��н������Y/@ҥ:ȅ�7��>_x��(��1+�#ýS1�4���ra�b^~��Gϙ��n�ch"-�H	��)fUsC|qY�?�k��� �,�E?�����\'^��d����X���$�K�����h>��$�1���L�Z
`��,�L�K8��;X�8�!��MP=�����@r�n�L���Cv|MD2�G?0)(m8ܤ���N5�)�^S*M}V������_w�a����Zڲ��ԅ�)�Vz~���Z𰘦Ab&�G��F�īi� �=�l���蠕�'C��=�����Qǈ�
�к�)"��iء��7�+���NC���*��
�sq�!�=���!�����"�-�6�X��'/��6����2!;�"La��{ ���d\{�b%m_�[����9)�?B�S��'e�����߱����x�vi`�Gm�\��ƃ<gaT�Q"	�O,gЛmjʁ����CƟ�3� c��zSm��`_(14��յ�E�VZ̬�X��n�b�?K�a���G�=��'��w&����=��g��-��~7� �^�B�S�����-1�c1t���bu��Bb?E�����7����D����y	4�>u��[C,��߸F�+L�����܄Dmі7�a�|��y�{�s6O���C��<65tZ&U�pEC ��R�`�ǟ�4�C�??��徛�F����^2�U�>�=T	�&����`�p�4�Y�^1�-�ȟ=���T
0���q���0�\s�B��Ҡ�0W6F� {�Bp��R:L�@k�������m�,���:�ADgg�A�PW���XW!�nXMw
�UI��k�PFM��ҧsɵ���I�1��t����\�Ί�X�!�K����>�w�|��Pk7��ܳ�a9CA�
,9~����G���[V"�T�/�!�rn��9J,?j��@���r7�F�u�0�V獐aU@%b��@�H�ן��I�^�'��Jo�<<�'��aw�`\��׽2����E!�5*��6�[Ő�R���J ��/�Ǔl�Kd�	��o��L������&�>%d���1HM� 4�se]Iy�H�^#a� ����n��d}s���MJ?���,ڻ�;]tؠ}�����G�p�h&_�ȉ��_���p����<Z@��K]�3Hb��[���	�ԭo}Z!���)Z!%��� �辀c�J�N��b-��jPޜ��">���Feߪy1Vٿ��潯Z�?��#��+��tv}�p�k\~��6�:8�(�ل�=	/�T���)�ˮjoE�i����	��s�eze�v!�C2�Z�o
�4 �j!d��c����;���?5�Y��#'1��<��U�� �B�%w7��zV�c�=������Q�}1����qn�p�!� ���;֞s���Ɇ�ΠB�1_�ׄ�ǟ�tO`�x'������<�(�E'����k{���k�+��q6p�Ya�'8܉\�����`ngѮ�v�p�����G�*�e�����=���_��X4�T,49k���J�#���!�3Y����
�}3���R��y�Mg�e�(>ɹ��N�ĦsT-�ޅ���Ȅ!�.1�xn@�.O�'i��K	��JXp�]@�D�����è @��[[�ζX5��ɳ�%E@�/{�6�ԏ�_���B�c�Gj����2��n�X��]�>9�J��H��c����>�OO�9,.���mEy��:� `z�2FI�Ơ���Q�y#%�䌿RY@	qA�t�S�E`�0x,G��x���'��I}�(4Rfﱨ/���U��f��A	�'�v���ǽ�X<��z���ʲe��s;�cek.���ST�8c�e�$�?6E�����Ĭ�q@��Z׷}��~<�̿�V8m����G�.2�D֊�.���g�z��0�5߂~�U~ut�83*ԑ���T7
PX�{�?�|�i�m=�O����7�&���4��*`�d��{.����&#W��Ǣ����$�pH�'\�"Bv3'�����A�� �zLC�������n��$	/�}B�6)K�����Cϡh�T���ٞ3�X-�:�0�C���I��)�C\�+b�����b=WZu���E^ޕ�RxV��]���k���ٗ»�v���>��qӍ,Ϩ�����f�����KV�@��:���8ݸQ�a�z6MӼ��<��C����8��ϕ�Jٔ�����%be9 �QE�[�,9��8�!�F���#^F�I?�G!��Y�u�=���]�4����2�����|���߶��@��kq��1�A��j��ܳZ��ו�4g8$��G��RR����a�BX������!U�=�44K������oƛ?�oN�c��ޖ��ή�X�j䝛ϛ�$�~�,���3uq_���>�Yڎ��UDٍ>2�j=�"�=��gD���)�ُ�A7��z5D�	#EJayƙM15��L���u_sݿ�v&��2�ƪx�&��0�9@���Fyt8���;�7�'�h�<G�^���i��������Ͼ6?~�g�QD0��:n�'9�[��C&@`�X��F��ǧ�|���pn�6���.p�٫��!b��6�Ɖ�Q��og�++�1_1��Tr}��9�N�� �ǃ�����;�&�~nm�dyg���&#&���W���j���c�`N���V3KbN[�V���S�N�mj3�9F��BTa��g����oqj~#{�1���q2$쇀z-9��I}i�NDb�;qN>z/N��9��=ܶ�dVũP����m����S�>�����ƀ�֡Fx@ݵ���v�)]RXx��9��d�`_�1�=��h*�J5�m���C��rщ�&"�c��3�;��ST�֞ݱ5.��\�	���
կ���`��d���X��Ԭ�g�U �8�z�K�3�<�)�1�dQ�ݿ��{o[L���f�q5`J�b���W�7$&�^�!`5�=�0�Ój2�;�������Z�ܾ���+4��xI�f��O���w�5ߩ�22'�Pi�'���ƹ������&#&D�P�!!]�Wf��Q�M�n!Y$�"R�NGJ��� ���>9@�ppɝ�z�������2E����ְ:�,���3�:GR�QN�G��[���B���:,#̸G	^`��D?��������b�^�ˈ>y>+p@ü�i;�/v�od?W*Ŵ�6��Fm�k7&Da����~��Q�}��a<�W�l"6��):߈�S�@�cM�N�ǻKA[e��Mw�B��݉mZI����3i�3˻�����Ik���W"�c�`CX�C�Ke��A���t��P�p8E��=/�h�ʋ�U�fI�\�-��<�v�
	_�#Q64p�$k��?�ItI��s"S�\���q �|�nb/����hc��ڷ*�)X�n\��yU�w��1W��8�ۗ����ҫvl���T��k����� ^K!H:���V�kܑ�9d���c.���%�O�:U�/���'�0UdrG�:�/���!�ܐ�0�=9O��Qv� pO�5���P#��I��H�xSMGeH����e:�9�����yHY�6���>u��F�}����a�t�I�Ew����)��`S'���d�۾���`A�0C�H�:��Z��,������*RA��L;�6f�ir�mT5�Zac�g��{���;��!sI̠͙R��6��հ�K��k�ŧ��w����NR����O�=�6u���h�X�V���0�t�*�#Vo��F�ms��u����n�wm8�ǖ�.ۢ��m-���~ߵ�^��+*�1O�������I�0ELL� Q�=26��wB�}�`dƜ���g�؄g��򜳼\5'+�Y�R�`�~�ڦ�l���sӥ|���."^�w��є}���ӕ[#2t��ی��X%T�/6n����|�I���h���ˌ�[����Bt�j.��K�%�)�:�E��1Lfa0���!Pw��{P�r`m���O}��uf��j�tЦ�}kA>���t�9�^���#%�h,ٵR��&ѩ�\el�|����VH�{w[�R��?Ŀ0!��=�ƙ�?��qy�#&�@�mR�L��8m��)�"^�.�a�}.�(��iD�$�,ɜ*Y:���h���i�mf�� S�ڧ �w]���Һ� �x������q�7�`F���?�/�9]5��D\�kr�O��������2Z D��g�S�����r~�Q��|�}t���T���T���]�k������'��^B�0h�{���W��K�A�/.M�:&��7�����e�_c�����6��(�|jv�i5�.���*���i%�LHi�w��ՀU_l�+�C�f�����K��h[��qr�/	�[�R��|x�b٭�d�P�K�"��lx�	Ӯ_z�o�$C�;|�=1g���ۡ������lߟ�Z|i��a��G����M�Y���^BIr���2�'Vn������`�\�v��\er;6C��'�f/�_oT-����%�`uyy��/¬˻|�@��ɼ:<au�YOh<�dv�x56Z7''�j�ziȩH5M��;��
�瞈��&0E<��Y���Z/�XVLۄ��C��3潰
�7�}{�:#:��S/����	y�{q�KU��#>��˻2�\��+�M`����k�[84�Ҍ<U�}�32Jw]�>~��~h�Jx�G��mZ��;���ƸirƉ���7��keM ?fR�:��J��g-Ĝਕ�Knv��]Y��7�E[E��F�좖d����h�흙ǲQli~	��"�9�c���y ��*�	%k����J�zJU�ܮ�'	&q��I27���	��rugV���XX�(Vr7�@��i\Jo|o��r��r���k�K��G�ྒྷ��ѰY�}��*�GɟS$M-#��a4Q�չ��N�e�
?�q�)�8��)4�4{�}ج'�z��=� �e�9#�}|��BwVYܻSfF��R�<��i!����㳀ڽ���"	��:��If�=���~O��Nv�������Y2���,n��O}���Tƈ�O��������r���Hh��9lo;���F{ߦk%f�×2����	��J���?wmGj�]��X�ܠ��q�1�F��2�NHC��hE�l�;�`G	�o�%l9�������������� ���9M4s�ɞS]���=>3EU��ӷ��7<�ا�9b���Y�N�T�I�.�R�k��8�d�lk�l
ONB��,'s�&��$\V��X!���K2�Ð �[ߝ�e��m���H5�\�}�������|F�t������$6����W}!+T��]�Yc�FG[*-���Ԉ-�B�{n$��i�X%�Dc������'�{>���׻�ʻ늖j~�3�{x�WA�b�j�8���OC�6��K�:������QT*@nN}�i/2]��"����|p��"�:VZЉ�9�쓽I:�$6!;G�� C(��	M+��1suR��ӫ�Ԯ�r#f8���l%�y�gy1mV��x0���w{K����<>��JI���(��
���ѣ���|�f.�q��'����.�s�����q�׆��r��8!.q�.�OGm������Tܫ�ݓ���x�Q�NH�'��u�HX�S�3��$�-�hE@�83>�'[�����!�}��`�A��TM7b�?�a��&��
 �vTI�({t<�3��7UC�V.*������`�˛#�!@H�v��ҋ�ɥl�ç\̚?�"�8�_�_��"m�+��%�MV�
��T�d�x������e���te����Hl�{"�'�[����TL���X�C������+N���|m��f+A�d��+�DM�	&/��fS�C���k��߫�t������r�a��K��[�!;`]oT"�h��Ψ*�d5Ǘ�OVC9I'���fm䡼g�Oۗ�Tt]����l@#�p�բ	��`K�^ ���'O8��`�;/
}@g��R�o	�DL���s�_�>k���\�[-��K���W�N
�r�B�e��(ѫr�B���5�R�=rM. ӎd�ۚZ����'(yF4���h��x~�ju�t�ڬ-�ܽv���o(�g�1ũOY�L��`��G.��{p�]FeF�7鑻@;���
2|�S>�1���.���?y����0��Ġ���1���X�Ǌ�$�D�ڍ.�Ȅ�z�:�óyM�"{��fn�-.�ĂU<֤��g!�U�:Y���Kg�1_Z�nyOj��(,p�\0�:�8
C��i��k4��+��|�%���V��Y����_C���`*&��;tU=����>}[ڊeI��#�KHP\��<��<����6��h�S�!�eo�"Lu��n�ѸswI� �"�	"��P�ՄCʒ�s��!�"y���TA�!OD��7���S���0=?�M�>��"��̏�Sgt�/�w4l��咁���RW��bX�t���c*[��p9���+v.��X� Η6`�қC�w�b�i�l����D)�7It��;<*�v�l�ؽ�ɉ�~��9�P�]�"�|-� {X�G����~]�N�PU��8n�s��r����I��MJZ<j᳊�S��-ַ��f
�����I�����G�¢(|ew�"SA9_�14�m�Xœ�����1E �
H�=}�7�/sӠ͉Ϋ��n1��p��G)���z
Vf�MÇ6�{���G��j��7�"��Ӯu>�T�Y��0O�6��^U�������L�v{�O�}BՁ�Y��|n %wB3�����u��7����6';_;��E�E��y7��cT���(�~��C��	d�c[���i��ʘd��_˷>�S��G��?���a�2v>t�P�D;h��F.TB�G��!�4���-��W��V�Aq	��؉,��u)̅���ϳ�U<{�vgiڱ�'����o�qe�p�_if>����� ��S�c4�=�X1A�G��'�������!
�9�|�z� a��#;�Ο�6�2#�a���p͠*ο�4|���i��0S?:4�A���ō�]9��]tB0��f�<��EAö��h�j�\�����u|�D����Gw��:�6���v���ҡ&����$_'v�
��
��FĮ��0�u�J����J��d�sA[`��7� ��,��KB%�T�s�BU.x�!��՝&.�����EΤ�+��ǰS�7�U(8�A�i��VTY��A��WA8a>��S�iz��������3�ܕ��1k�񓸷�#V�T��L� ��`'ȕ��R�9�|f�3���bA�Z�Q!#l�'�!r��h4��33�<��fS�P�!�VuΉD�ׯF�t��E �F�Uu��/��[�f!���B�����$����;�Di!��ߒi���;�y�+wY��K�=�(��d�^��/Uf#p����4�/R��JE�/�}m6����i�Y�[�.y��D�V����׊����Z��P�'*�Mf-Qd4�("g�;x��l`Ab�x�4>-ʀ�g��p�l�$��H?u��J��ȁy+��5Wl�����\��� ��&�"u���ϣh�A_�%`��S�\�@��黺������~����>ͩ亨���/|@>�w�k��݈��3��
�\�Ȁ|d֣���Z��M�̓��Æ�Ts4��]zE�!�'�r���%�8ك���^�]+���4�l�N+��0/�l� {�S��!��M"&�s�����Oȏx,�2O�**8�?h�
�(lׅ}*�d�;VYιt��%��,K9B�|�u�b�}�4�f�E�8B�ӑ��T���3�ȼ)NƯ,��c�B�ĦxGJ	G�D$��g*��uV>]>N�:^���M5��
2���B����曫���_�T
���M�N�Y(Oj ǁ	�w6Ɛ@	[qI�������$tF�Y����'>��

7��8 ��~��#���6�bQ�����EV�Pׂ̎�3�^z��Q��U���������cPޢS��?�G�f���	N�58�4�!t���ԯ��7�D�!�7�^�7�Ƞ
X��3e��Ę��s�t��ZH�����;�rl��ߏc�27������{�e�nO ^q:b(�Y��{G���6[=�\���V�[��S����~�Fn|�`E Q1.�!�J\jX�z����-}�&��nU��G��/l�e�:��j;w���z�MND&�<ZL�l��q�z��"��}�M�[_4�ʑqS%T�����w���W��~?N�8==��j�#���Hm6�E�x*{��O�04�%D�>�F�0��H88Jp�J)�)C�����5��cNK(s_ �������yޢ�G���K�"w5��]��05��
gI����ỏS0F���$i��cx���r:�rp�|���,�:�:	���C�r!.)�g-�G��@Gc�,,�W��ps��Z����!ͤzy�����w������P|
/���Ю:���x���д ��`�hL��!���6E"H�XK���2G��ȝ*N�"g��.dr l��|�׿'�u�y*;��x]��ѓ��x́��i�n�'P��� fg��!ře\��xK15��ů9�ʸ|�-��<�[���b·�<��#��
��2�ry�Ҁ�B�*}���(���/=�VMR����Z6��Y��F����U��gC���wُB��j�l*8S���N;7�=M>�/D�l�z��,�����|r'�L��"�ޔ�m{%�O�v�
�0`N���Ν9�5-��O���Fh.�=�9�h���x���Ԋ��?����hd�hvMڑS\ޗ��@\��Gb�I�B��7��?����5���(4��wT��z?=��m[�
o�1CVި�S�"w�ge4�2�`e>�aaI�OيhY0`N��$�e��'���Ƌ�?�e��^%� �2PeA��J��).��N���o�4���4l�0��J�+}}���d�������gny0�qKS�U���>�N���D��K�t{~�ſ�}�&�±H����WB��_��)�g$���Y��?��҃��C	��� i<�Ԏhi�G���1W6���G��d��;����T��:�Ox�pE��T�-�,5�5(o2���?��=�\'1;�>=��F�3B&5�6T$��K܉FSKb���N�u�49�G巵����|Z7x0��=�c��B��x'y�g˚:.�]�&J2I&Tl��:F��|�D��L��?ҹ�e�HqY�Z����Vpa!�DE��F�+��.
�s,)	��Y� w�M��-�st���	L^�%�K%��N �¥K����a���e�A7eV�+�	M�.Z:� ���9�M��U�o�,���*&��
#-�h��Y@[��s7�zy-�E�=eVl�U�fI���z� !�����1�7w%`G8F��/�)���(g�=��OaՓp�P��}�ل ��ur@�U���.�IIPg�&<]5�(TN�R���y�������|{BȞv)O3	�O��s����1�
�ʴ{:�LK:�`�ٴ2�#E ؎1��n;�P?	�a-�g��,{��M�":_uz�6#��f`7�ȭx�!q��u�[N��V�������8$z<�#�������rChE��{�Y�9����|����t~W�SٱF�U����+��� ���~مq�b�̓=k��&S���'p YU��R��eJ4U��]�l1X3�(:�{V�x�{o�N˧��эA��o)ZRS;��X���PQ;�P��z�$���*��$Hu���薙��> �����h	�=��Ɵg%���&���Y�'Wp��y���nTu�2�/�����c.��W]�� �e��e�]
��_I+9q��y���&q���h*

�Q<:H<7�X�>�[>�-��LG�(\�MYbƵB*�/E4��д�oR��HML
Pl�\-��:�uT�Pp�#b���]ۣqe���{SꝐ�Y������t�`A�U粫^|{J؛�g�}��u������6� w�|�Y�� ���4�G�Mk�N$�8���#b�Pr�ǲ��U�Q�&�S� �k��)Ť߇��L�_ '��/�q��:\C3A���`bi�������Ƣ��g�S�}�P����{���x��yb��QNd��kCǦn�&	�~�.��?�Ӹ]��WRZ�Щ���t�~Ϛ�S.�*��d�z(��d.L��$֯�JmcM���%v�B%H#y�#���ϝp[V]��@d���ު�*�2y�����%
�
؊���2Ty�*�,z>��	�\���ʕ�h=Ҋ���A?s�P+@a��XJ��q�Âd�$ՙ��D0e^a�D�Hb��p�����C�Dت�������p����+|PS�����Ru5��&�fj���{ޏt�(�*�#M��T;�T.������?^������ǎ�˵�	J<�*���N���9\K��5|�Cf`mوmh��i4*���~��ZB�Vw�B�3���T%�=IR����,�CTsf��~$b�Z;�@x�c��u�8���>�?��؃������{�P|(����.�;��#�n�*�Bh��=�a\V�����$�N}4�țW�x#ZJ��$����(�X�˽��D}�v;ŧ�Y;�I�Д\ۋ��"�����7$rZ�u�:����f�6djv��V^�!�>Ayy�����ٙ ��(��(�i����a������1�f���?�@����N�D�^G��$:mr?I��T��h"J[K%�}Y�@�l�����k"f�ie��̚��$����|ֽ��d��s*� �{����Y�=HLAõ�+��ӡr0;"�`d�_��r�1R�H�����_Z��re �$�ს99�g��?�T�o���2�{1t��h�1ԍ<��yR�f�]:�'ly���}�YE׼����v��鐝�ԕ
�������~[��3�(�I�gNs��c�q9H6�S���\1n�T� �tu���,v�~E:��WA9�U���,�oG��z�	|;��\���	Oc�o:��B�<ڢW�z���P-�����I��=�Jd�,�ܱuLZm)K�k�C1�>����~Yz@�����,�
\��ƚjNJ$�T#ﵺr������>f���HN^T��c����]�#*N�N+��0cI�Z
8v,�F�K���X�ظn�G^'��Z_I�Er8D}1���<י�AW��[�w���A�ON���Uz���N �\����J�ӥ��[C��Ptc�,�eN�2�-}����4�x��ḏ��侺�U�"0�_���q��-���yʴ�G��7<ځ����Q����(�Q�(�����b��'7�C��%`;wP�=��d�3y�R�����V�1<3yFwN����1kz�x�(�]lf"g�AK�EN|Z��('T�Ђ����������~w����E��7�	����g�I���n}�me�F��by����6�{	�`����(��NǛj�i%3W�9�8�]o/{7�DM�(��9�%��hY'>5�,���޿
�$U�!���R�fU��3�H�7���u7�h17z9�^�i�9Vj���<ɔ'/z>ɼ,ଟ=F����R�!cb\���"�LR�'�b�Ł�{����,�3=��X,ʟ����h�z����	���cq�l@��.^�1F�'6r�d�����X�r�K9F7n��OYL�FL!�\����U����#>qT��J�+vR?[z�%�S�:?�{u-eG��C*�>[$]+��G��v&庭����vT��ڰ߹�Z�c�Z �YB��'ċbJw1g1B��^�1�M�ۿ|^�sXZ-�j4�h�⮣!���$�����(�����v|��,���>+)�Vw(�,J<��O���J������}���B� 4�aE��;{s��rk8��;Ck^N;4t�U؏}��$v0=�x;����V�Ha2bS�#0,%oז7�jK_�b"Gb�X�*BNU��$��,-d�t�)��sAo�[�:3�ct��/��r-��P3��w+K[+����������&Y�ʯ���S)5y��pނ������{ D��#^��Q.%�I4�먕�^�`�6{�������]A j��E�S��"��]4#%2`;���U|�
̞"�r�� .[F~>��W֚_��	���-���)��ƕj4ImL)(K�/��(U8��������u�+DcP�]���~#Scqz�
����n�'pH|�&ؘ���`䫄������p��1ߡFIPCh�<�֝�k��@P'#�����6����nv�eFG��9�%.�ո���6�}�!|��8d�N�v0�F��bk�u�YJ�2�!��܌�p�UK�&V�8رY��W1n���1{�Vsg�Ӣ%Re��#����=��1��Qx�W�Y��m+�Wt��.Y�G�˯��p�T�$@� h ��$��{�*�`�ٽ��lU���`��v��;�Tp3Se�ȑsM���G@?^��5֢az�L�ef����������r����k��(���f$S3%��Qُ�t��"b��O��eć'��'��9o
�<T4WAH�P}�Lg%Ņ�E�Ȝ�� �}Th�< 5�.��u`�<���oz?�l&���Q��NUa���`��U�M��#K���H�YQ�r���J,�|������CH�\�|���f�ů���u��ʔ��#-w�7��q�Bt�.x�n��E�~����7�'��Rb4�6�$ŗ���4�R����LP[�5����j��3dyP���)pÈ�4���4@��vV}�����E����p�hiw�� �w]�1v�=�W!,և���8�/���:y��Fc����oҠ�\~fСI��[Y��0���*���H>��f��F^�ެ��b�Ms_����d\ �;�Cc�ݜ�y3�m�y?���TO8eQ�c&�ɸ��/Eͤ_�R6+v������l�b1����,���}w�6b�#�5,F��qD،I�x�Y( z�q{Cf����[�½F�3�������e4���k#���T�!?�~�j��Bh	FT��hH�O!��=�����A�l@�t2������2ad�BH�@�7,R,��i�V%�Z#��;n�RM��>XX�A�����~�erj=��B��=�n)�$\KZ�%$�7-��\�S&S��F�u��U���טc�9S���-~\]m���Ĵ¯����jbƴ�M�b�?Gtra�@4�F������ӕD��hM�~AtkN;l�)�_�{ �<f憎�z�
\*�_�����I�?q��~ V)�܂uuY�6Dg(F�%s|��`����;���D����v'�����y#�X��Ī���qRꁡ�l�FIUrp���X�%���)'Ɠ���X��Ɖ*� !���`QdD������{�%�����Bc���A��Z��O�_<�M�>>���K��+A��V@�h�+�,i�h�)+�Yd(Y� ���Q�7|�#���d[/�<�!.o��XV�����=!H�Y���e����X.�9+K���ak�o����/lt(��]s���m�H:8~���M�r�;ui���I�*$������^�n��2Q��rٌ0�/#B@�`Ҵp�z���(�̛������)��մQ�G�E��<��įe8L͵����e��:�{_ARt��o2a�r3�/0���I���P�U5#J��C�y��a��n�
5�=x�	M.v�#z)~����m}L�Xux#4���P)���?A���e}������_�^�,ȳ�ۨ���&|G(J#�qy�Q�I�b|S����B�L4�q ��@���l�n�n=OW-�t�k,��\��(���d�U�A0��� ��~$xBX *^{�-�Ɓ�R�2Y����i��i;��'H����\�E�g��y�l:1E1! l��Fd�U����p�r��R�����G�?~�ake�ar
�{p�9}�A~��;R��|ϫl��FVڬ���lo��A5]9���a�B��&����r�y��*ۓlᘶg�ï�1���m ��|Ա����Ih�_�U���x�#�D�\��v�tA����}����&7�:�"�sP�B��R각�KN��M�8�*�_��&�����u�#��gvn����-z�?z'�W+�z�p��+��q�}\�{f���{��u�0(�G�z���B�X͘Kz)�2��w�xZ�]F��QD��9��]��L85�8�i����j��RsOaP�Xe�06�n%�+bya��G���e����3ą^I+7�D(�An���	�b\�jTJ�>5�oI���!d�P��嗏�P�w�vʝZ��b���ZK�@�(r�'(f�7�dtݑ�Ȳ�f?d��4�
�OI��Y�V�yוB5C��9����;qT!:&��0 �=X^zTG!ʲ��(T��\ �H*Zݭ��o%E��
x��[@j
�,`}���/���0��D�vKĺ&�k��)�M(h®c��$��5�At�`��)���kOsE��P��%�cp9e�e�t,=��GL�h�PZ�>ٳ�ߓA�b�S��G�΀���:?QTR�NK��tPܹR�+`���p�\�P���-]<�$��)~~HJ��ȏy��iz4]��g}���e+Q\��n|o�+Q�O��\��tg\�ϴmP���9R	]���&�R�mn��סP^��{�Yޅ/�uf�X�e��y۝�r(u+�-ϙm�����WJ�������k(�Uʹ���@M��H��K�4�������,U�5v;	$
�FT��ZE�_�b���1�����0uY~��+�4\�|~d�F� s?��W�3P�n�^��K<���� �u%BSB�(�8WL7�Ț�}Q�>X˼�~RĄ�w�-{�N�'��5KH3����尃؁�t�wd	|0�F�ћ�$�!���Ƭ¯>�pW�觃]F���\�Ø��f��Q�G����	5>�VPe�ʐᨺ����gх\�[�	�ѝ��rИ�:�$�$���΄%�;c	�����BH����|�~5��#��l���Z�� vn\'S��y�L��D2�yƳ��f�i"�5o�`��2jt��x�����T���C�:���� ���&F4����4lֱ�"��4|��2�W#��������B��E�Լ�B��9�� �Sp�BRO��R���\Z#���P�����SBxS6�^?�OE�����Z�G��ڐ�P����b���hU�k]�cW3��G�akԓ�2Z�����m�����t��ްA\{sm���� 
?���;R!⊟�����j!�G��/k7N��Ò2��-�K��і��8��d����p��d~�~{�f��p}�(����%@�������՛�� �Y���dic��F0�h�)2���(�dw��1�~"q#-A��1{�`=��e�8Ƌ�Ŷ1 i�~�h�BMN�P1�M��5�١�7!fqB���S�îB^ 	�u����z�ፈ�<��E�>�M�u�x\.�BAH#�t��d�p��K6v�v�u^)2�R�6\��1#�̐"������^W�/c.Ǘ(`%z"���~}=��=u[�Z7�](�܊�;��͔�#K
/���,S�F��u�ȩ�����i`>�2V�e����8΍��3,���C.27�u����7K9�6�ٕ#�Ő��V}����ݎ�����
�8�����>ځ3��?:߯u��,dg����.Al��v2lw	��A�b���&��/��h�9�0��@(���R]N�m��2f"i��z��?��s�W^g���H����1Ҕ�8��{KM7ж1ɞk�fy\�]��vs���АFt 3�������<6��~�b3��q���s�2�Eh��Go.���_�Ė[Џ[O��h���#_P�s�R��Q��)�m��؞���B��, #����D�92�Q��4F��!	�wΫ�1�`Y�A���I赚�9O��D�~|䄕�=��xqq^/o���6<v�K�qh��!�O�B���̒53�zFVm��J�2E���J�=ׁp �-�����S�YY+ؔaVa�z���}���(�=:X��}��Ԏ�T�)�+��6�m����e�vmiQAG���ePO=1��d�M�$�ykaN.��F?J��&Ir'�F�`N<օ�[y����J�DB;�&�����$�*:���e��H��!At�9�7a:�k��YV���ÿ�A�	��(F9~�e_��Hz:����)y/O�Ȕ�(3>kI^���L>E��l�#�/^\�	 a��/,���YR{�?#ٻ�sH#!}�Xy���K��DKb<N�Poa4J��S7����8�YD��ҫ)̫��@Wv���]f,b�Um�p c�Q�{��*�S��y�U$x��<�aM۱(� @f����Lk���e�%�O���m�e�_��f�}���#E?�5ٹ�(�M\�����6�d���1�~�����z?}��Q�#�?A�N\�B������2<@dvv*�+�K�Ǳ3��e_�y�ZZ��u�Q;5BR�%���b,�'".���igȶ�x맾��PV���uΊ��b]4��'��<��4I~��Xk#��\��Ju��Å�{�$��&��i~�6�3��~���G-T��M�6]�i�'�j��/ ���Դ
.�`{R�Q_Y�J����2��j��s/|���/tp))�|��98��-D
Juީ��<�آ�֚�.W�=��M���E%1�3ҫ��"�P�B5�SO�d������������&��$'�Î����ڥL�DlK/7�=l|V�͸F��F�o�	�
4���h��/	��19--LyQ�C0�l�����30��#�_^^�rr@����]�Q��#<rN��xS�BGJ�}�oPQ}��Ӟ���K0�FS	N^����.nrnb�oǞ�� 
�%��|��40��V��71f�p�R��%p�q#���o�Z��S��W����+���7�]��v-o�N��$]ո0#4��ũ&�9��!�%�����d$����ظ
'���;�Jn ���E��>4�"���kO�/� �i�����'we��K~!rX�9i ������M�i�_S��̌+ݺ䷴ℙ��,x��"�g<���o	� }��$�F���!|�}1s����b�؈?��}w,"���s�QJ�SXҊP�*eT��"����D���]��{������2���\�á�D0�n��ypf�K'ϱPX�|���%��M�W�v:4��u�N諤3w��I�䟏W4����k�ԟ�O���H���U������Ͼ�E�Z/��{�J��wF�0`�%�oI�.��
��Do��>Tf�E�M�/����h�`XG@Ľs��O�I�I���;�,탺���?E7]4����Z��dO��3����}Ud���G�w�,@��-^�W�ް�tH��K�����J_cs� X�(�f�"�����+������k��)w���W��mYm��J�� ��<?v���۵$��"hB���kx���b���\vS�U� r+�+��<bS-4?�)��-��B\ke�K<������R�>pW��[�Q7#��&|�"*D���3�$ yp�2������IC[wAS��5��:{X�z�3'�t�i�u9��Dl�i/W�I��21F3��ܱ�d��:�\L�V�^j1*$R�ǚ ��'>�W��`dN�4$�g��I��\��-_��^�W��-�?�i�h���%ʩp2Dʹ�?@�_��c/��`
U��x�Q���)V�FG�D61q��\)�����[z��j����(�۴#�k{vV�=�}o������=%��ѳ����[��g�t�Nd����$?�6� �e&y�`��d	1	���zF�٭3l��P��#��5�;|���eV�+=dͷ3�v��G�H �/����D�aѵ�b�n ��� ��O'��7�;�L�.���dy㯊����}05������2HA���lr�G�Ⱦ@�ڍ/$H��t�(��~ʑ�N�l�[�q�͒��a�)e`���>=�3��ӭ���3)�J�!}�.�(�W�T6��I$��8��D�(H�!b��dO���*�H�]n���!�u�AO���������@!º��34)r�ub][Æp~p���͘t�Y;�z"E����͔z���;��?��L4h/E%���-�ni�j��v��ݠ�u���.��tpY��t�<��R*��7�o��-� ����f���iZ��8��y�^�R�Ӥ��m|{������P�v���j2��;���g�iC�X3��,��v%���y8��^௃(�-[��'/�8%���\-j�q���ͻ��q��tT��l[LoҼ[�PĐ��ź�A؂ #�(���6M/S����e�����i-���27{8���Ai��$2�t�Z�����vu(m>��0l>����� �n�$\�	քB���B$tN�˅��n~��"�ir8Ԫ�ᔘ{	o\��T	��l\P���f�'�kCc�|�$�{Q !�y%!wAL���eOb�����f�+{�V���Q�Kb��M�`b�D����;!A,#���hDO��m"%ɦ��P�
"Q�ԤJ��$���\�q�W̈́����A5��𿯾ro�p�q��3����v��ki��ڥ���{�A*`�X��_A����KYt��#u�I�1�� Fiq�"lC]n��w�fܫ��� �%���#h��d��#�L~eo��	�Py&9S����*���=����U�P�.�u�u�Z��u���k:��c0��c@�P�pz�W�ġTGEP�j�y���E��L�Qy��LOeM��v��wj�U��4d*i�YE��W�$�3�RZځ�vw�[W���5Bm,	��4��������V�'
�{L�?3�������+ڰD�3�sI�B�l��<+�y�F+#{TpF���#��V��R<�$�x���<�v�S�S-�ω~������/0h������<���<���7������gг����opUl�4�aX�ki�xd �? RGZ��j�X�ȃNJq�(H�� �����֙(^���6K`!}�`LS�9R:�s�Z˿ãc�h� ���M�z�WC�Z��q�$6rNoJ��:����])0呎��L��C$n��������h�1G6�(�r�#�sUǟ�|?�'�JݵX��f���b�}l\��I={�!�j[t�>��8�(".G͐"���-�C�m���B���k�#	��T�w�(`Xlʓgon�fB�6D����Df�C$��by�T�%���s��|u�� F$��OP�W8S�SA�?X��Œ^|s���N	>B�Q�єW�J��G�\��QR?��3.�T]�Og����K���ҧ�ő�^�K�6��x
�+S%�QB淟�
�	Hz��g�Y������\v�8�61���3�����h#nA#jf7�l�[��Gֶ����27�^xp��w��S�DS�!얀s2$tN�.j��T���o���W�s�^�'��N�b{
�JvM��t6|q=j駒���Kh���`����Kj�dKT�a�����`��O���V��)�'�7+�7K��(b�t��zj��r����l긏~�<Z˵}� ��γp$�'.�!�P��Q����֝cc���Q�P��ք*߇8k���׆�����=�m�;�ը��3�$�i����x¥+�cs��&�?-���]�����knt��?�;ݝ<@��`�wu��<����0w������({�����������
O7�:@�G�<�0�MX�'lkwa�z3��\
~Vx��Y�*�,$NZ�b�:��G��~k��M3�h[�d΋�'8t.�F��������2�F���5�~�Ltً�/8[������g_\��	RlP!c/��Æ�t���B��8r{�G��NŐ��d��Wc$w����qLM�F�����9c&o�D'B��;��;��2�3�p�A����<�'�v�E���fn/u��� &�������87�$-��(O݇B�ޫ/��֊��-X�--����36 J�΂��";.5&P1�w�����U�ܖqq�PV�@(v���#��wx�F�5�2�4�g��"�͟�i��Z����4�2I����j���D-B1��� �����.{K�ƾ�<`��]���ŵ�n��3�~���a]Ms3 k�:P�H�T�],j���$�mN����d�ql8���ԉ��tj=>e&(|�Q:[��5L,e�|+G�I<�K�%@�4/D?��FC�0�&S���Qm�L�#��f�{� �T�{a`����7���"%�M�\���F�s�u�B"q�42\'Jp��)�Τa���&S/X�	_�Vk����8���?,�Q�\��Ztf�EG.��[b�O����t���f��?�g�4z~�&�ݨbG̮�W��h�ߝ���R���!	5�Li�ͫNF}��ؓ*eIe.P�B��$McK�v`�#��ۇ~�����3n�DT�� ;5�{|�Bճ���s�H6���i �U�I3BZ�\��k��˙�IK�q�b���-ԈZl�)���p��=���K�uB$�c̋�sP�!D��=]��X���(UlY��~�g]yo١�ߝCf%�Q6�˝n^���pvKT�R *҈�P��$�����+�~�A����}-?�4�+��_��f��<�g�YN	Р3d*�I�ͧ܀���NH�ܣ�߻�fd�����a9�r5���� 9N�S��`EȀ�� ]���=���a��چI�Èen
��f�,-EnK�/7�z�{�Ӌ@ub�Nq=�֟2���fC�|~Ũ+N![�s�����K��7��O�)���7ix����M2�w-�F�S�+BY�]Ozw�#u��%6�Xn�ɾL�ދ$�#�N��!w�h˛��|�~�@�����g�o�خ���k�gŧ+�9�7�e:E�3���(l�	<��+~;<��s\$�.�{J�=C�^k�v�����SE�L^˧N�q�Љ~$���=��t�)qF����:R��YwT�q\"��ɍ�I�B��?�k� �~&ؓ�ވ�*.p� e�2�t6#�[��ʫV�Ӹ6��Nh6q k�z&-��&�{=��*XNoc����u-eN�u���FH����r;TpKw�_ ��:���:XJpXR�Z�W��3��H0��6��x�5e��ZJ�3�L"�|�)���k.�x�tL��w|8�1@��/��Y �o�C��5��X��*��F%�V������n�����{��M�_�>�<��S�ơ��Ns(���:დ3s��Z�5G�������ϴ��<S��5�7[0���T1����P^pW�wK�
 �����*gps��x/Y��+'f�$?g�]�`�
�^3�=��V R3p�܊��>eY�zӨ��е� ��'����7��:Z����n���e�)m���Os�F44�/K\ 5��V��n:���'��*r|���'�@�h�l�P���o]���h���*m��y�t։���xk'[����P���Q��Jl��6U�|l?��`��b@��.R�:_@��&;�9X�+o.��VaQ���wb���V�=@Dcu�����&�İ�n�B�m�t�V����y͐]El�0L��ɨ�i�⿝lxb�K��U�8KP/�.R�Y�Bv,fW��|���n�7�DXù�T�4yr�=�vQuSz�
K��G��9�S`�
r�Q}u��^�{�HW;}��Ⱦ�;�~��=P7S�0�#���5��5�i4�*m�S�0嫕Û�4���J9����+�X��G��e�J���K�"�K��Y圍�}y�8E1��뚐Vw���s�.�e㊡�KI��������`�)6��F�N��dn-ߙ�M)f'+6w!!�9��$%�%����N�5Xb�9�z��K�^&��06<9گγ�F���)�ڽk's�Xn�x.N�$ޗs��~V��S6��u�į���}m��J~���޹�}�m��5��l�Lr�X��C0k�^j_B�`���fE��ɟ��{�F��&�ou	��xkS�	��
���A.�e��d�Ƃ5��	��PŹϽ`�xV)v �+%Ju�4��g��3^ny�aA�O�LP�>�?I��5LS�zA%(���}b�^1t���|��*���z���(�.�+�zWȔ[�\�x�8��)M4�]�Ж�m���k�V�X"W'�YspYaJ���e^��.��D=gA�|m�W
I�P��i&l�߅{���қ��#j�+�^���C��+�?ƛ���X2l��B(85���L�d��ɣ�**��(etB�³dk�PMI��6_?��1F�ދR�}��)�2�R_0w��J-F��g��=	w�\5!ܴ�(�E�(�,��|@V]mN�:�d�2���n��M�ۥI ���&�L{��A�&����| E��|��P7���!2}���#)��o��ї��;�ζMh�>Ӌ��N_x��s,p��!���|��"a$��B���(��2d�E��Ba�%/����z*ؚ�;�Čx��>�SD��ħҾsh[W��H���N�UB� �2ī}vx׷X>���M�.w�<�Ȝ^���:sG�/����`�T|7�N�7���f夦���6PwaO�S���,A���Vi��T
Ֆ�=4�V=K<��XZ �%a�Հ�PΣ<8zz⯢���{`F��5�������S��
k������t����fYO�+��ƹ���6~��azz�-���&W;"�So5{��|�}������W�:���,l��������@��d�n�T��r�`s �u��^��!k�2j30sr&�\p�XF��R�~K�[�W��ɑ��
Ԭ�#��_֪uE���2�>����w��=�W(�ԍ0��"�c�ʾNç����XN��u׈���G�<jb�U>��.��.��;�jL��e,��GGmQ��,��2NbG^�M�� �Rg�~�>dWl�>��̀:fƩ�_�V���z�㓶v�@k��E�����b�������B�Zt�?��6�";y�1@�zp�\n읗�{��ڀ7�w2���� ҭ�D�n�qSE]XE�M6��l�����i	%I3��W�&�R����W�n\�j�	��ab+F�����j�]!*�iR �w�3���^�u	��ˑVO�<+��B�b#��m�+��n@���z��<i�7�UW:e������h�_��B��K^�ΏҲ��U��j���BV�������j3v63����׍=�EbxVX㒖��j�حCv�;��缉3�b�žRi�^�w�g>�3����y?}���� #{�ވ5
��.�T��@�G*_{��)���'HXF��N��rB��yd��q[K��0|�)�_o ����-�팷'v�i�`�h�g[���,��A�UG]YT-ؽ�`����F����w����Y<�#5\h���ҐO��3����ݪ�� Uy�'�W�\�ֶ6Mfz��>ڳDmG@a0�.8l���Y�Ol�S�ہ@���9�uo�^���wdc��.?�]�Y$a�5G��lK��Y ��5>0I%�v�U����0����|�P�J����9��d`Ϲ����[�,�{T`7��&��с߭ov\�|�����?r���:OI�U�sQl?!%-Ѩ�2>�I]�p��P�ҩB��ƥ�C/d��>*��l���jb^�_����'��ݨdV�.c	�Ҳ{�L�hc�r����U��;�hؕ�!aj������D���VƇ��;a���WdJж�ݓ)��-�ސwU���j�&�e�~X�L�C�ʈ�*:��,2��IPP��{޹"�O�^6ܙ���G��i�=
�;}|)��bM�K�X�]����l��탛y��T���`?��j�,�6Ƹ�f�U�q���&���#~� r# D�+<p~���3ӫafu�_u��c��d���J(���_/zC"�p����e���{Q?���D=��
�xT^4�3r`�x#�f����ʘ��/��l@hщf]ށ$��S³F��W��Cy�ݍ:un��52"S�v�m�*�����`I93��~Q�����֔�#PgTVmu��^:��>]kԙ.�`�[�g��x�v,y�pTk���zQ�S�/�^Yy*-�mI� ���z�����QbOb�ߠ :�|,���0qCq�+X� sP�,�����\��~��ݷs�����ĥF�/d�,�� )�+�Pڹ��R���7x��LF�A�(~�>!w�Ls"ɓ����mb!S�T��TXj�] e���ݍ	�:�`��[E�X�1:D��K|'�>�����:���M��n^L�,&��l���aɾ�ER
����	S���w����Z��E�vEǓҳ2 ��:N��0d�*!]B��99=U���/��)��tR�p�F�+J:��y+��5�x6���R��z������=�	�Ո��e�m�^����IGAO(�]�T4'X�Jㅕ�~Ƚ~���O�o����
���NƧ��QLl�Ϸ�?�����n��!�2��e��>c��4P�ms%AfJ7х���3�G��bB��>;�G�eOӧ��ݞѷ���xԅ"�����yC���	��Q^��;��ǂ�\���5�R�ؤ6s��q��T�����;z\���w�"���%�p�����
����=��.�ڥ�4Z������q��#����	2�	��k������<kL%va}���5dt��Pɲ6aD"���%jr+���������N� neRA�"����~A�-�䑛;����$�]�S8r\�+��]��f��T���i��EwQ'P�_�M�"l��0K��kr��#X��#�� ��0/��̏X�\~�ˢK��֥��\aޛ�xWK��b5��x���Ʒߠ�-W�.��$�1Hg��GqA2!Ot}���+���{��3竱�6��H�řny
�_��O�0p��l�M'$��@Kk�7u���&��u�cN!�����/�;|�w��4�DiŐ�B�MY�3/��:n��w����3�+�Zx{;�RsnL�U����[k�t��?bMߪ��z���K����S| �<,&�8|L���O�9����I����=�#�\����w�RSe%��p0/��	Uu�<��8.�T��b'��+f	s��gM}łI��>j�#/gA�K��24�vA�\�拮
̣�sEص�ݕ��#*�2W���Q%��s�f[�U2��6z�^B��Z>gj��셓�v�@hq����Mg����u�N����a�4.[� ��%�-B���쯕yRɩ���}Q�%�82Q�`}�n\�-�V�e����r7k�~�4�I����cZT�?6=F>B�5K�=͘^
�!!����3�:c��1�_JB�Ph�!��yUM��ְ�9��W�z��&$�M�����ຐ�`K��ץy%��`��4V)�1��UR/���<p4i�z� Ka���F�,펆PN��2{�G���=ų:�v�Mj�1�t��9�Dã�Ɣ3<(���[�vaŸ%�m�2%�7��)�B��~�����5�(�q&�)�(~*j���g�����p����6�G�4RvI�Ǧ%����pY�<	�����ũ_5UF�F�� �2K�.Pr�֊jP�j�Gq�Z*���Y��<���`I&��|d�̀[�VW�ҏ�(R��sȼ�Q.#���QY�бCsbװAǶ���,��38�|�9�E̸�&D�o�E�0[ʫ���S�}��o���bi(O �8�.�_G�@���Pg�L��Ǧ9��@�B�����3���͢�Z$��8kM��JN"� %wW�*ֿ��ԩ��Ox�QNrj ���jl)�Oߡ;BJ�?=�\P��5��z	G]\ri���~���Ǧ�2e�%G���J�WQ`h ����(�zz':N�tS$1&�<A*�d@`U
#t�r��EEM�S��L�(�rᅰߔ"����#��Jg�o�0���ic݉���=ic��X	�nB�����v�Ʌ,�N�.��0�ln�M����Ea�$c2ƃ�/��!�Y�*n����ÌAI�sH��B��eaniy]�p`u�UwQ1���ZL>]��������O0�^
V7S	�a�cƄ&��E~�~@T,��jwM}��N\
I,�X^���O ԍ ��b�'����k�܁L�<�x�����)��@�>��z��Nչ��soc��iDɍ4v�q=�]�!�iv���߷��L�$9(	��S��y��?���[�R����p �N0�kC����<Rn�lJo���iux,��n^i�]<l������)��Z.$y#���LBX_��+p��� jv��q����X��=n�h�n�*���磈^L�Z�/���<�|�~6.��
�#O��v�%�:K���׃%�e� K�f���`*SY�v��	V�hY�v�E�T-�5�7���R��G8'�d6u$1l���z�����Ġ���O+k��>��8�Ҳt���z��*�[�r�[
�(g]��$7�i{xcQr���j/.++6�q��S|�0��~�+��jZ�q'�T)�W�������b�g!Ӽ���k�
޳��r"W����Et�+��-HV�([��{߽�u�g�3��h}3E�����0��5������$Q��8ÉSwyq�}���K������V<��F�V��e?�ʕߙ���"䏉M��xωj2��V?ݳ 0�i��`���Ҡ.����V����C�k�GB+��)"�ٯ����Ν��l�"��EEÍN`7���4��H*��k��zY? �e\��E���T�*k1�g�C�*=l�L̓<��#��y2�&BB<�E�\�ȅ/�%z#B�A}�]7��l���}E�U�B�Y��h������؆t�DԱ������}a��I�"\�ܙf�ܲg ?18�N!A]�V��ɒ3�8�1��^�X���}�=�qnv��N�(�+�/�_y�^o�9��{�#����~�<J�����uIrN-��f��]���yhB�l�:����fY.��ؚ��|i���z�W���%�E0�MV�"C=�1nI�X���b]�2��ٹ�'z�.�i��T�t٨�)����"���	�H�����t��I�d% 2�ғG̗��:o�{u��ir�D?�d��p�o�!iΰQ�"6���Z �Z[4wH@��/�bFG�-^���|� m"�<��c��,3>�[}��5(��oR^��ao�y@��
�=���@��:�gؙ�;H��^I���t��K󰅰
ɼ��X�B��@��J���O�~�Il5tk�ƴF��o�湃N�cUOʫ��v��`1�)�g�"�FT�x�x"��<:� h?��62��$��N�겼]�
�@�����ӘY��u���&VӲ��&=hʢ�|���<r�u�/ѳV���0�5��0y&<
{��l�R�d���ʚ��g�v�V����)SG�z�Ov�� �J��d�,_@��kE�
(w�	=3=7��Ä]�|��]���vK ��1�dg)d�c��w���tF���sơ�W;$yBp���U2������y6J�R/�P��x�N@5��N���-��?�`��_���arq
�� �^�oa$n����~�*@���%j��SdnB��r�ěѸS���)���8�	{eq��;���O$���k�՛�7��Ujť��#R{���s�Vϲ�1����N.�SX�'��6�\TR<���&�� �?�������>���1���5յ����T�!a[T��C�� L�ɋ!�=�|	v˟$j[۰�7P���}�� �ʗ�'׋����͑޶0�!���1��p�-�f�Hg�ƾqЧ�7�3����e�C9��Kd��aG��P�7c�Q�K�����>���&S�#���n�Xnlh���u�O�ɰ�jkk�s�n[�^�h���.��{I�M�"G�/�f|�~z�
iM�
�n�2�� ���@���9��d(��)�4;�7���c_�hNJu�D�RlQ������_���>
G:�n_�i��Bkf!3�4�d�<�zBN�|���q���u!9�� /IX�#w�"l(�>%AҨBX84�"}f~)���o>�Y����9�V�le�WoOa��]�x�=J�29ƶ���E��9��)�1��|�*��PL*:�(�9�O���Y�V����[Pw7�[e`a�z]#	6�,%���ŭ������>��������0-��v
vx}?�R���rP�?�!&U�X�\�:X�>=啦��{�?+^E����!D
D���HIv�+p�P�3��ğ^�T��uB. �V�+�_�LU�1��S��C�N��b���]��j<��	�X�����"O��?�W�ފ(��mdܝ�|��a��*�o݋i�o�%~�׾���(���o�Y���@��Ģ,� 3� ��<��f2�EkiDQ��+଴�w��h�)D3Gp7I1�|_��X%t�oete�i���pq:�M_����'J��Ur��c��5�D��w�����ty�Gs7��B]# ݷYHR�Pxvb��O|fwO�7оX�I��RK�+�j8h�Ӷ��P�P�=_��S�|6,3x����+mx�S2�%s�Jۄ���Lh%s{Lf,��iڿ�\̆|�K�#�@�&>����*���\ �Z����;�� y6�=��"j�WaK�#&�^�sՈh�Ni�%*e����ٱ�=؏;\�:�3��&�\u��Զ����w���?t�g��x�s&�\�`~����(��|��	X�f��q2����Є�� R"�o���`�/�[G`D�khy+J�exv�`	�\��ਫ����G���,�N�Pztx'j�4O"4��H���W
����9�/�(����4T��O�/��9�!3srG�Q4V�*��f�H��e/4ǋ
]����x���I6(s�H�#S�YC��L#3YF��7�U�\�B���[/�ܝT��j0�O�Q��#jM�:�ϓ�m�Z��2�Δ����<��(w��V�+��j�ux��n�k`�Ca���m��8�RqЪ* 2��P0c΃G�`�P��_`��ۮ��GrO�1�t}\�,k_�άHRom%R���?��Yr�&neH8��c0�6n��b�Q�T�P�}f�ö�����b�;��+u�$V���ɝǅ�ʻI�G���"��NZ��.&��?��H��`��RO���r��Ӝ�Tu>�<6�SlY��P���4�C��� 
P��w����u%L�8��'T;D�ň=������֪8���c͹�i�;����1j~\2�y�M�A�w��(U1�T�<o=��c/BE��lT�_�h	����荾;�}uh��Pb�%z�D��8���<�af��I&|�Z��4�BN��.��x������p��_���^��V��Ԅ`\��A�	$�fi�E�!�]��)z��Oe� �������urlh��з�W�1��Il1	)�~ަ�ǵH��y�w	���B���.�����>;�OZr�'�q#4��<��D�'0��su�=�Ed98�Zv�ڦF�<�V�r�B�r�i����ʢ؊?��#E dVO`��g��F1��T��Վ�
Ϋ�U:�^�r����<�Zvm`�`GJ��Ģ
�������v���u�Y e#��� �9�8��h���������&�ٿ�:��X<�2b��OY8�q�J�m��=�RW�4�\�\��q���];���mf=N_%�"-����WtB��8b	u˗�1�!=�H���F�E��C����I]�渚b3 pfG#�vx5rfU�����a!��!�\R�ԧ�V�IU��P�5�
,�@}�V��/�Ӄ�]�J8�m�N���kiMc��%|��nľ�}�{'��W���n*�>�dy��1�uyqVVI*	3s��5��q;2w5࿱BM��<G�������I���7�w���Z�%1{|�����d҃G���Im�D��WW%�ώ��6]+}p{�%M��Nԅ�Wk�k7 n��pp��^�ϴɥ1���Z�:�av�����X0qS'����i�+��У�)%�l��r8�$%�v�g�3�f�,瓥ƭry<�Sc�""߈�̇���J�cKA�<�b�����"-%� ��i�~�Վ�g�^��b�Z��x���w�D��d��Ѵ5&ILL"?�� Uw�0�M����}!���y~�?�%y��DB;}��yPUk��4F��Ϳ>q�=F
�F���q��l@��>Y���)��f-2��.��cX<�F�p�Y>���we��&����۰� �4�{�7��L~΀ĺC���7@);�+��~����E�����Q{�!�1�)�lp��ɀ��Pٯ��Ư�|�����AŔ�d�&��$_��HxICaث
��xV�����e��yV�3sP�x�]������j W<�G��z���N!��`��-'/��r
�x��y.�[�'�6�8�#Y�,q���W*֌��ly���uf@4]>�J��#�q
 �=0,J�yƥ](�Ϡ�����bb�v�����|�nx�;��p;���<�"�?�i5P��F��� J :����� ����
b0�]]��OP(���.�kv�	���� �^�dH�@�AT�'v���~HnyE����b�)�?��P�.���sr>N��C���8�/�L�Ub�?.�8�|F����i���CVi/�1�v��uDu�j	��-~�����4鉤�]��o4n���J���@�,�ailD�_
�[s��w|&	y�,�O2(�aۊGs�K�W)֗��u��G�A5;��Q"���4�G��
�N|=�<����A��/1��TS]�I\�����3�OU}��S��{����o���3][Y�Ð�K���!��) �M�� 7�u�]Hݦ{פ���ޚ��͒c!�$�a0	z���x���Wu���#�v;b,"����B�>n���bV��	*��i��.��~bC������1qJ�p��^�F�.ד,,���P¬���4��R����>�S���k�
�^<ߞ;G�~�5_{
�Qw��*�P���/5��uW{��rPR@�\�T��r#���0Wﲼ�{nڻ�v��G��b�R���2���&ľ�vc@�59T�XoXܰ8W4��a���ݗ�=�]���q�hN`r�f�/T�pZ��0��9��(�S蜏�+��u}�K�l���X��|&n[r|�	��n��fQ�+�_0O�l]��ᘩő����	͒��
oى�L\T(�UB�|A�b���n�2��*��.�mS�87�|�_A���5���c��َ%%�{��6��|v��X|�w�b޾�1t����4hU���M<�>r��ʅ���a��r�{��r��4q*������'��93��6�(U���'��>�~��Ex������d��kcBf*�p��H2{���P
'���IQUA�Y#� f�hԭ��d��K�2��ъ����gHp<!j�IvR�ˋ=��*���(媶�X� �s���"�k��<U�h��Xi����&WK:�������Z��1sr�+l=��ˮo��өX��9�T��u0���ɱx[ʝ�w Oշ��	sLr�t����d� �x�\n�y��*��tTP�����޿����!��A�Qp����v�4�Y؏	4r��e���S�a#|�a.U@[�J�B��=�����3���۠֒M;���X ����$������nl���>�����3�WR9�~`o�v��Հ9��\�2_�;~��;e�R���-`n�<;\��u
ǯ��l����?"[H��������[`�S�G��+��*���D�U�� �O�}�P�� -1���^ѡ���J9>��5ol�@�G#Gy+h���^9S����Ch��غ���#%`��@�������ٴH-��� %.%.u�Ɓ�'�҆���B��(^2b��A|��`H#�t�&���Lu,��r�9s �=�l�e�V8�.�+�rK'03�"q.��i^����t�
B�tO&靟\�-�X6��(�/1�'��S	w,���r=c� ���L��>�$��j�~Ͼ4're���Y_!~�	nh0��h.���5a=�fԇ�VX ����Ł0��$��6#�7wb��Ô���c� ^IK��D�>�vW3�?L��E���XiYK�������g�U���sS�vB?��syR�")�D�s����2fR�$����;����<ã����㬭,�gAQ�����H!��/I�� T��iWґ=Bă̱�x)7ܱ{M�����*!iU�XjZX��/�^�	w�8`rBz�q�����;>>	p�Y���͐�䳧�p���M���Tw����2�� ��H���].�ѓ��굇$�p*��w�kk[���$���o7'��ڲ6,�M�n�%v��x�!��ӽ�����X������w}�FE���m�c6�j�>�ǹ(��%�l2����2��c�����bn,ÙH$ߊ�ٷ�H@ܟx�lHC׏9���ga&К�����n[Ԓ.�0�ފHJ��b�3l���G�7�}��K��I�n������$��D���������{��f� (a�
l�3A#�ܦx�R�u�7���E]�Lg��/�%���܀�#κ_�R6�g�U��qP%R�M��B2�(
']U��?�H4Sx�Vx3���R����U���Iv�f(_�3
So���Y-��5�AVR).�e�<�d���b=��������F��7P&>%�p�l;�8}d?e�6sGL�)H���|ɘ�7'@�]���$B`+�뾇bRim���R����j�K�G�����LK x^�`����M���+�ď�O�5���):��GR�<I�F���9�_��g�22p�K�"�g��t���iB��C�XA
<��us�gp��+�mn�u�\R7�I�bRRz"�D�q���d��J��\0�� �d	������,,h�y�|W
����>Z�2�4�����s�UE�L��S2�Ir*p��M�)�|*:�}���{��m*�9���.�[��5Pݝ>�1��.�9$�����_�&'��yCN�	�6�=�P�5��˝a�Vb��E�D��H^�1�ޑsćLb�d��g��˩��`���ճ<�/x�x�.�&�[ʬ])W�7ny��RxH���i][;<��"|��鬺��*�V���1=����,X�۔� �u���e*�z��G����N��[X�H�Hi�l���q�UT=�����ӆ��.�1o���Z��g2��h���]|�4#��E��Z�!��:�2�l�J˿&,�6m7�P��7��Z��\�/�i�U���({Ř#?���T֣c���T�M���6�6��� �?�����Dex}ٜ�P�=�v�lt���1����2��0��P(����Q(���|g�v_!����=�f�]"Y���^1�?��%�}�rg�8]���58";�����!B���%76�� ���ZH�rw?$���z^�X�Rq�����<5�+�6�� �Z0�| F�̭��KI�%�|�5��6dDC�TՇq9;��R&�B1�z�SMkAV�*��[޼7t���(��vU�e� ��*��~��.4ᇌ�GF�jC�a��9�I�8�a{�`�zA�ALJ'�b��v�gVY�i��AԆ��ip�a@j�� �qp�A.��l�SH�l�.Y���%/�C_���t�:;d�H��m��&­ W�k^��ae�4���6r��sI�S�iß��XL�O��nIP�]-f�(��w��~j�}�c���F�W?�W.�g�_��VV�(��K�qgi�*%K�������EU������1���OY�Ծy��!TU$��eU�T�'�$_�7��k���$�G��UmPƳ߫��.�<�_���%�F6I	�S#j�Ltl�,"����m�9
��Ҫ1�y�0��0MGb�/�g_�F�����1�$�J�O����Ԓ�@��S𶞴t�{��E<����������@dd['FE�M��7`�h���V�55���(7�xM.�x�nCc3Y��@{HA�R�R#�ך�!�N�Ok��3�^R��<����M��è(2�0e�5�	@��ґm�i	Ѣ���^��	��W͖����� �/ ���w���bTF�V�;��`kI�^K��,VMн�����V�-Kg��f�L�JW���A��A������?S��*Nh���լ¥kMDgX
jp�P���2E����t��ǒ�s��E6:���+��Rs���tr�@x%\���V�Z6!�e��C%cq�i"���ԥ��L׫>-����rcô��bv�K�͂�jJ�`�Kз.�{'��_L�̘i5a�s�S�*7��gb�ж�y"����U��k�����i�H�4��,������Jr��ҕ�c�e�w�}��8�%f+!�>E� z�������\���u�YnfK!�/x����U���GN��h�q�b㤟�3��5�)0*]�������Z��?vy8qŚ���np��E8��o|-����o,R�qK����@bT�S�M��¢YAګ���[����*`�1ZAA|�(k1���TJg\-�!���t@?\_��r��uX�ͻ��f�+&�st*R^H�K �ͻ��Uj>�i�_�.:�L�������u_�J�e��[��ݒ!�^7���t��-���g_W��Ly^��A��q$׾>CO��{�x�1َ$�����h�espl��p����Y���u%c�[qD[�-n�1�g)��{*��]"G���}"q�����fŔ�A��ߠG�۶[���8O��<�rPtS�\�`э}Ɍ�ʻj���u�Ө�+de���f3�7�~S��`�'cq_���Lpj���<�~�ǷI_����Y�D�+Ō@��Tu�[����,�A��J�^� �y+ʉL�Ē�-��QӒ���`�d�m�\��x�i/Μ���ŷ��|uV>/'�zb9��~���S_�������y�6�l�o�P5�k�ub�C����?2v�3�ǵ7����T٪Iu�<�������F�Z�i�����b-�0���?ܖ��Y�>	��O�>v6�CX2�:��I�1.@Jd��W�%����-�C�@DY������l<��Ò�Z}Sm�L�o�4{�h�?A� �ŷ��B7�(4�v�"$�N_e�|�ٮb���04�˧�Bm�󚾖��~.?�!~%�ح��a[!�U4�ټ"���13WR�iMd�y<%����짦�k��-YN>|uV*dzA+��x���<���^Br�j����[(���nݵ����R����\�)�����2M����·k+��;$��2P�:����z"�������X5�hIYcM˅c�Ďn��GG�a��q�T5%r�����Y�c�:�=�2��G#�X��h�&`�e�V3z@�oЎ�^���}��F#U������a���[d�fA�my�W���u��i>Һ ݅�9�=h���P1.:��w �&�?�$��uOo�kJ,b�
�E7���"/smYF�;����T;D³��Md�5��זA�j��өO�����ȉ�gԬC9�ّ�6c
��n�0��qO�L�אD9|D����%4��eDqu��Z��reSL�,��+{craq�4"M��m�*��?��G�X��3�L�y��M��&���2��D($"z���`R�6�Q&��[ �9#�w�>Z�^��{j�Z��>)aP��8��h�PFj�˲�����_���>D؟����f�Ƌ^��ݏ�q����rA`�i'��Ǟ0��$���4/�ǙD�Q�����r���x�	ӣ��;)v�;�T���)��a��0i!I��&#��z1P��L�;a�%�
1���I��rK�9�Έ�8s�x���5���NJ�a�'b0�y�)t�Bی�r�O�7�LaIu'T	�Cr�er��
%���H��E�H>��z?݈_K�{Af��A��L�/�T����I�
�(��$�e���E��q�Z�cW��ӛF{�sBu��=����M\c�NRZ
���C���ǼS��6+ߚ�/�6��v	��dv}���"���B��-b��co���<(�A|���$��qY��9�q,��aY�Q0�#�Q1������+6�=�~q�p=҅�����2R�F�K�#�>�;ļӸy�7�V���t��K�cS���Z+�3,-ƫ�5�K�Y�c�����C�䵽gn�p�?2,���A<<�q>D�<>A�[��cT�f������(� ^ږNj�z��8�g�g�yU���>�g�f��7�~f����a�l&�)de~�f���#���ͭ<C�&(*U��S�ؾ>��Ƣq��������8��z��h�|4�E���G]���ݐ��z�2h�Ʊe*Ni�}5+��+l��ts�2��!�-%j��E�T��S'��b}�*�V'������\NVk��&�0d<���A��+�`d�M�:�1�aN�X5��;�m0���,򯽂^qH|�[���a\��,P�`_����z�����`D���aae|� ���O����ӔN����Nզ�[�˂jzT��ҝ���3���ZI�^ꢤ`S3�c���-��K^0���]3��Yh%E�h���������c�d�T6���3�m�]�|Z2���C}�@�.�fDn�޷��f���RW ��s�|JAK)�������!����9��+���:�-���>˂7\��\(�I�б�,+w���ĭ���6x��m�Dr�f(Mֱ--�r6��t_C�����'�'Rfg�����%ٔ7ǖ�ҩ��h�w7v��(�2xX�w�Q����&�v�F�rĥ�"��(�V|��$_c�;�W�3u{���g��Mǉ7E�������wU&8e������D���������p��yx9Tk���9�f��Q��[ (e%A/�a�T�F�g\t.N��,y�0�vr��4��KM�8o�|��+�-�_ �+�Z�/PETQ���
��1��ዽv��BԬk�	�Y��i���p?�Q���=�I����.�W� �a���M��J�Y&��gPFߧ0T d����A$�
�/���N�VFh�(�Z��,"��2�R�Y�h���-*�ʁ4d��u	�z�TW@E�{��f��F�Cę
f�d��K/�s�Mw����>�ӨOMP����jP̲��tu�(s���&�K�7����l��ۆ��_.{���8�k��ݯ��Yq�3�2q�wn�DԵ��z7I῞mU�]hr,:w����'c�9i���V������2)p|-|ε���d�34�S}z�~�/5�~`���0Sz���eܪ���'�V E;��SP9�'�d���=�]��I�.uZa�Dw��<c�lȓ.��;�%tҎc?�N��.i+6K�F�爰љ]|&���� ���a�XE�Uhg�����E ��oCoӺ���Y_�	��@��̄����ĵe�J�8�
[�,R@u�P��ds��@�>����~y{�Z�،��7m�3��U�Fif�=B������W���8���Y�.����6AW�O��\��L^��{�4�N��RT���\�oX��w+�j*�hˠ�q02�hY�A\���������|Y,iUGu���[b����̸���P1m�-9_��/��2�7c���|��-^5�/����ȣ,_�[��H���E���y��1ݎ晾�#����̌�n-VYW�JF|%����̛:y�l��-^�@ ��2����~��~W.z�Ty�uR��Ϭ�;���/�d��T��������1��R��5f��~ڝ>���sS�f�
 �4o�u�c�����e�@�v̓��׀�ʣ��S�T������`EI���V�x�u���l��B3(���ԉ�4`0�.o��*���NS����()om�w&�1������m�Q�y�k��B�ᯓ��<a�C(�/��6� � _�
CMhE)6E�p�H�JG����|� �LP��g�)ݿ�_�� x��Tn=p���ț��F\�qP=h��	aV?���3����qqA����OԺ#�����5�MZ'p$��Q����]�c�W�����Z�j�]�l-`[_m,GIT&��~-n2P��g����}�w9�J�����
N*2��.�TIe'/++�J�a�\"%1�`��u��J��뤞|j}R���o���`|6��yOx�?��{�Ɨ�&�]
!L)Ͱ���x<��0KlJ�U���o|�b��3��<Ѐ���4���}'`�]m��z�-o��� sB�A�gh��#%;q�_Tu���Lֳ���/d�	�MD�?�?�F1�5�Fٲg�ifJ�K8��A��)ٲ }i���p.���o�W♒Kop��7���%6%����(/��5�'�k�>~�aU��G��]�r�����}6��m���&��}8��i�[?ќ��R��w\S�������s���M$����H��*�b�H�\*���0��$M�����,]�7�����{��E�pƮ �� �8�u؉�!��'62��߭ s{$V�؂�o�ǆ���ܮ+_++PkU�� ����5��w���)ek���A���b�As�))/�㰠%���Z��(,6�6#�yQ� �9�Z��*� E��wݟ�r��A���{϶���1�)RZ7��Tfg��{p\ż&L"��45�C��!�vi��X����K^(�������+�y|%3������
vh�5b{G[nX��s��S���w����&�jr����N;oM��Q�Kz���hJ���q/!�S�F��/����IQ��h3���k�r�N���0[,[�2,�\��G@���;��\�!����ۼ��^$�d5�W�Nl�9�K��˫7���A|�(�A��ƃU�9{�d���vL>�����yd`LH֞�q_O��ܤE����H��P��K�e�Ām^7���l̔U+���ˑv��m��VR�����[j�V(�{r$S:�٥�Bq.3���?�<��+��i��9"5�I=~��[�`]E�^'<���AЛ����C�`�x�L��z֝,0BG��/�.���ke?s����}��z�G,A;&�5�8�n�n�5c� ��<Ku(iDF1�ֹ�;x��Kq��� �[�����GFXb83���hz�����w�*^ =d�b���ڭ+U�]�
�� V�#���,��Z0�%��>��sһ�4�pT)� iYrW(�`A��brC��%y8�aBlR���AHX5���"���ȫr2,n6B�:X g7 �z���t�3zY��]Hk��p��\��+�֤Z�V/�2n�.��y� ��ԫ-���'/M������s�Ӵ�2�*�R���g�5��M��f�w�Φ#�����?N-��]*�vKw��,H!Y8aD��w�u�B5f�N�!+�8�p9f��bw6�bo��wF���р�m��r�k�2^<O�m~Ӑ5���͠���ݛ��BC�%�����°I(��3q8�����CZ+����z����|��"k/^�C;j�:D�
R�<I��@�����<����8(�&��Z�1H��˻�R�3��56a��*ఓ�*��F��e!X��`�[,�X&~7�����F���0UM㇋G˸[�����3ސ��Sv������F�n������;֓yU�5x7�����O�����4Gc�*C����p��Z�vTPcr,��,`�]�~x��=0�)�+��ZH��m$|a�Jq�o��U�2{�>�r�$e��>��.v����1��W1~�jV+�y�ș�F'�I�'����m��!�]��<�L�Pv��c���`�.�9d �^_U��^�2TE������(iT����5����_�����28l���wt��uy'FN$��1ƺO�)��ْ�YKش���m��2q���5$��0����1�L��:�n��B�X(>YK���c��Fad�/���f?c�)LDM���2���A�6�����,%�J��4�L�Ŀ��-����P���6B��H��C�gn�@��1=�`��]���g��Z��[U�@);��1I�%)N�55�Go�H������"����u�2E&yK� �_� &M�Z&��	�)Ȍ��	�g�
��n�R&%����;�G�𒚐R� D�|�����oP��<�A���Ӫ~r�~z�JM�MA��V\�6 �G�Y�;'��C�VZ.�R���u~^���M3��&_	z��}��w�"�]zt�ݶl!��S�K6=�P�T��C�vi����3��e��8��t#��1�ɳ�S(jko �nO�������~�c&V�m�벳��67Rߩ>*����Ǔ>Q�	? ]�1��\6��X�M�I�u�������]$������z��*��W�ư�����p��x�u�j����NEɮp��Fp/�T+.�1��[,��1��A��!���5AaZ%ߘ�[t�slM��]f������V͆���= +����M��fU�E���%jS�&��?��0g`Wឦ:���p�w8�"[.�pcp�[�͓�;S{�L�������G��)j��<��k�R�B2d�(�»l�>���E��u��5�!F1������������I�m�3�_��v0����;�E���!^�m)6fOeH����bi�8a��MZ` ��Če1��G��?I����t2��;�x,���	��R�*Ą7'��*<������JqE��R]5�]����2�������l>���4T_�{q9��!���Inn'	=��VB�n��i����v󮑰�_�q��&LY�ͥiqc��q��gU��<��� ��δtc�2�Lw�]�P�)�=�'�91z�+-1kqy��a��Za6���.���ّ]ʨ�����$V�O��~��b��J��g0�"�Q�A7b<&��{����U���"R���;��2CG<푭�Z�P"�7��F�՜<��A"��z���H�pf�����H�w#7�����Fa��GdC��m��~��F�\*x8Se�hz��sl?;�t6�M����ɂw|�4h�H� -� �6�<K�]���a���0����D��"�U�ZL��˸��@���2����=���[ђ�vh�!8��ԑZN�%��%A��`gD\�X�R�o�n�ԟ�e<�}6� �wgȲ��@�,��g���+y?Ϩ�M�h
�h�B�qAke�Ol'���E�h
�+�����V!���_}��~�kC��:7�=��D�������u�R!����ˉ��H�|1s��T�:�����|ڰӅ�����(�`��h���Dp��Z�k\�wNs��Sec�(�����N)������ �ŦEl�ҽ�(6��ݳߢܛ��{u�Е����?�ɻCr��f���w�p�I��� J�q2L�F��F��Ȫ����2�A�We�P,$�Q����+�����{8��tƁ��d����՝�hjΡe�.���d�)t�f���%�����0YDl�Y%��7ِ�1�!~i"�����"�=�g�Y��Q�n�tD��
��%�M�FɃ�/�&a��1������)��b���;{?B5��Y:�B���I΃����s@.gF���a8_ʘ&��i�z��*�+�����u<�c�Ƞ�>�Ť����).�B!�w����/�`J��������Sb��g���>�܃:T�z'�ֈR�ALBo�y����طB��	H��\���=���vŻ�xv�����2�63bq���,�f0������ܼ���-�+�z�>е����e��>mi���1�y�	Tgr/��-�d�L���k*T	�-\�X)���h�wQ��E��E�w�Zh�Fpi9�q�L���aLWl�� ��n�,��N��O->�����oE�R�@l~hP�ń����f����O�q�3�����P���vVc�=����k�gO˛H�?n�u��mP&#�g�9�B9�T�c�^4؋$5*��T��!C������$��~��tY�~Y����V8��ľ�aE&�^^l
�L4�qʨ�|y�f"���dk���$�V�!�ՖR���P��hx�cc���g#�Y��ɓ{{�V�(��z�b^X���E�s� ��*�m쉣����tیvc�L��b��&�R��L��-&6� coYj�\�lU�$����زv�3�뗩/��4`�,��W��꿦{�8?�C-�:�ZUq�4���n��4P����},����_׃�m����"[�}`�Mv*�TDLF9�ã������9NU�#�|)^�s��N���_���MϹ��q��!��i4'����{6������x+�lPٞ�o�����bO�t��|Y��Ax?��ʤUv�8J�F��}�a�xA��Q:U�W�]�%��7�$#�	\����ߔ��49�% S5�ЬHקs�p�y#]U���u�A�?9�6�0�|F.��潳i�~J�V�|l;�h�Q��»��v����8��?�o�o^��3C&h$Ȁ����	���H�q_-:%8fS����?��;,�C�^�)�[�����S���Q���^[��󙝳��$[���/*i��|�XO�t��R��������^ɺg�i��i��M��/������Q<�*��Sڃ(�2p��:m�@q�3�ՙ���o'�	��nQmˡ�\O�q<5���B�?�:Zwk`7=j鍥b�Xʐ:�.B��O*�݌	���y�[��t\'�&�j�����٬l���jD�>I�L,����` ����&��t�1�[7��ޥE��k��Pz3W���A�.{S9On{��W¼�Q�.=U��g�6qN�����R�a�p���ܘ�Ug�Ц�ʍZ���_���{'����+���]u�*�wHh�)�8��t��c�v�gwD���3{�H�z$,#.���&��H{+G*bY�.@BMT����$!F���yz\&@��C�𪚎����@�D����
�|9�J�f!�@�-�4SnCy.v�J��(Ďĳ����hވ�ܦ��!��A��Ar]�D��ʮ@��6��Դ��%v�}>�`7�n@�/t�+������Z�����Tq+z���+n"�sL��O��&�qX%܁�q'<�n���K�XcS�����cߟ�\����޷�&.'���E�u��}�ȶ�h��V�l�oh���r �pA	�X��<<�(M����S�7�r�i�:��.}�� 5ԏ��A>�}�����[r���{��hP?���\�iy�)�I�D��2k����Da�4}�HB!墷�vz#
��Sj����=�<!�����+X-�����
;���m���]%�xwa�'�V�b&�-���y:�������@����g��;�����lcB~<J���G�5��]>��_��y�Yݨ�b3Tf{��b3`�뵞���d	9�L�4c��C�m� �˦+Q��"������Z�c�s.�O���8�"�s7`ؒvȗ� �CV(*2���ٹ�-�?+	B�㯓�`Ғ�yq��Z�}���P�X3�S*��/Ou��;��D�~���=ro���gF��O_�����n�g����5Ѐ�N��h$ w
����@[N�}�:�d�暇C��(�0h�E,9��D�v�A�5�RnK'i�瑜|�����%�H#��2�uJ��ȿ�+�"���\�tm�K������|)�r����|���hƸ��t�x== �����ks�
��r�E�A��4+鿡ܰ�����i-�e�Ʌ��fIʹ�;�^��xc�E��u���\Bn�UG����U��Z���N�J�v�}��L�'Z��6���9��6^7S	.�a.H��}�[K`����8��,gQ3����2��� �k'՚�&�V/#�M���wAnN�}0��P��[G``Vq?�1��d~a��@�U��>�jw��}��@%�#,��s>M]į�t�Y1��WϺ84V�խ��B�v�u�E�ܞ蓬����<ɶ�Ӈ��g�[_�3��A�=���+?^&j���l'6����x��|1�ت�w��냅�<��B�E�R��������	ǯ�A�i�o�!�H9pDG���-V�� I7E�7���-��@�=�Fݎ9'�]���6ֈ��G���?�x`�RtM芥:�A�R�4���Ӫ����Ek�@�$} &�,��q) ��ᭊ�E���४�l��!��	|��d�@yc�Epx
�l��N�l��X[����R��q�Bb�fA?6u�.���t��8�cWk���';%H�ih���P �(|����L%�+�����d��4�hc*u_������\�?D�>$��������^LB��EҮޑ]�����P�J|F7���n�V�K����_M�N�ޓ�D�y�;K ��'>�y��b����L��<A�e����Ϯ3C=�&7^q�G|���O�ϭW��v_��uӒ���X�G���EĒ��1I�O-�O���F��(�v�����TENo�/��*	ه�i�8%�:�
�Յ�U/�ј�ȵޅ?Oe��f.�c��[i�:��������N�I�a�U����3�ߐZD��Gf6b�`I���w2������j����+��s���8,s�Eo�sT����N"�;���Ko�B�_a���M�[��!�2�Γ_�[(���ݓ#��er��7X.��đ�������q}u(�nʧ8B'�����-c�W�P���D0!Nm�l��b�{�k�+�@�+Q��=	�b��k[�
Vo�V��y$��(��4�`�^�QJ��B�~g:+�[�v�m)n��o�����_�n�b�U����w�L�2�C���O@m�D�x���~�|'5 s��r}h0dO�D��E�F�т��'_3���'R��I�
[4}��/���XU�m΃��q�g�j��F�?�Nb�:+��}��KI�~4{�|��'9+6�F�ߵ�W]-C�G��F���&S��݅���x kR(:=�������(�]��V�8�x+l�Pت����ӄ�_��6
�b~�3�#w�v�F\[��|c��5"�@����l"�J�gߒ����"µ�X�O��ţ�A�;��'�e�3�a����q3��y%<��>�J^R�\@'�	F�Q���{Sj��Z��j����4"^�gUw�q��T]�+�c��	̂"��H��&���~���o��e��u�������[V��[�� �Ꙗ���� 9>ɩb7��+e���4!�ߜ����=����x�sy'�[x�v���*�l۪�g
���MQי�BMl�`k�	V��_���xw!{�R��c�#��@Ğ�nԟ���Mu�BO`1&�*���&���f�[z��汒u3PK�5��Ҹ٩U�i5Ϯ��-FK(��f�0���] �o��-ד���;�Uۈ���06q/^���\
����	*.�ɖ(��?�^�jEZ���2��N��!��@'�ˎC�]���<����א�g@�j�Gy,e2�_-P�1h@v*��p/���"�Q��ߛ��94�ڇ��~��_�cX2��ʤ0��G�g�h�k�UT�����6-|�~�� )'��c��Qo�y/�).�S5{qk����w�ȨC|��>j2Թ�����p*܆@k��v�Y�ll���a�`D�8��iN��G��~���q�o{}���
� �)����S_�,W����ͦ"�"��Uv��Z]���=���a7�<�8��*�:3��M��kQ�:+EĭG��� K|�N���^vW>7����f�RӘM/;�1��;�5(SN�R�݃Bd7vT.|��*2�g[޶r�u'�Y�񮽦��,��̖e���j'��6�.���_1"�Sku9x�:h���j�4��ǉo��^�ԑ�����*뺋�7���[�����[��K��M`Nj̼�Tjs���o%y�"�UF��K+t�O0�V�������}�ڋY�I��|��T<�sHa'g�Xs�/��ު�.
�c�Bp�Q�L�p��x)E����E��J��w'ʫ0!����H{��?O�ࠩ/��Z�c-�f�L����5^.	�Ir9�j�i�>Y>}���_R�F�f��z�3���ߍ!�:���E=X0�<�W�4���`���;�r�ɣ�G<�O{�o^�w�P�e�\���mD�����Z�*�USuŁ1#t�wv.b�<<��g�}�6�-�h� {�|��Up���J{�z�v�D�L�lz��6ϒ�d�1�9rW� 4=9WNu\�AF����1����w�#���2�|�����2�x�#ǐ1�e*��c���ބ�}��A��L.lqM �J�kN�\�Q��c��HS��o1(�fi3���YUܛ!��5`,��r�V�M��3����H��B���x$�xl�ݸ��[���oh���$�.�e2�o���L6e��I��U������D܃���n4$�-L~C�E���k�X�k�Xty�â���{ }ڷ�����n�1�[]#�B��5ol-���QQ��$�#_�@�-"m��2�+�4�53���2]��dƫ������hq����W������5mK���g�kPc7�FӉJ�s�)�����:�Vbg�VtG�Xz�	Vt�r	K�܁����a�CY9��p�ϟBc�����7$.~���;�vdi�}^LJ0~S\���&�|��Bf�@��������U�>��v��^�n�u���ª����/#��z(�q4�fp��m��͵���0�L�J�ۓ�N5s��kѼ�xA4e�?T�c\,7�Q�ߧ�� ��Y;m�ْ�_��bE_U�������en2���q)�N�&{�뽇�l��"�;�ĳu1F�e#�A6�ǭ��Y]t�C����Pb��u�v�nb���W��gr�hB�:�Z�h�W$~�����k�}Q�o"Fe)i?�P�x���83���~�o5�ݒ�.��A1¬p/I��>�06�!��T�&���~�(�����ͻ�sr�1K�~j�_s%�G�Ba 虓σ���0� �س��D�*p��\��|�N�-��Y��`���A���ؚ�)A9��F����sd1gwcj+� ��h���ȳ�zGb\��N]�s@�*6��ſ�Y� J�f6�)��t���̰��FG/'�;-�Xv�t7�&C�5F��W�{���4@\�y���3�4�Yc���<I3�S���4c�4u"��=�[V�TZ���5*w���Q8j�ȃޞ��3L�F��E�A�) �����y��B�wվR��)'�9�\��K%2�{M���a�9�切���:tYf�����O��86�375T��е1Qm^��Yy����Ƨ,A�0����9O��kY]$U��kj�Ϻ�ǣ6h���Ǝ/���-*Jϕo�a< ߸\��[`h��D��Ιf`�=�	Z�q�W���g(���V�@�����.����Q��%�e�峡 �Ix�xjߖ���u9�!p�E��b2bAq~~�5�B�+.�w��0�u1G�v~�
�jt� �2��&�23���L��W���@�k�pfޗ�*��A^�������P��̷�n�x.��>ؑ_f0�(�~�������lG��җ�"r��P����L���?��[G":z?�/d�#���u}�ʳ'�~4d�$�w�~�n�P(�ju��c�(��t<ͩX�z�O%����`� �L��b���g8k�G��:X<@���R�[�'f���,1��WGX��\��|<P��5�ג��ڥ��을�#���O;̦�����vcC<t��z/�r�x�� ���Ά�?�� �JgS���\|��t7[)��e�`��g�wp��K�i]@2;�w�>�d�x� (�I�[.gVMh�bx��O�H�%���7�]$[ӺB�����OJ_�>z�$�Ӄ|A7p�ɽLΫ����jz��z�r�L�N{qr��Y

7�jǁ��]7����;@>ro�i }�Q���N]�ͷ����9#lgvhH����RDp��@���" �ɝtzȅɟ6�Q�+9i��O�^j����(3�Z��&�o�p�j:�oF��<�k��������;���N��,� ӱ�F��l�3����!�dD^rC���{�+��v���ā������{�35��2�l��3jŕ�Ϭ
�&��"�F^Q�TՉ�)�kÿ�g��\æx�c�#���@b<�i��Jy���G�pF�\�&��Z�x/�/�������wuE�r ��,Q/@���:�3B{ߖ~��9��J�k��#/�:S:��Tk��&w�f�-5�n{����<l��L���V���؊�\���Z�>�/�N�Id��g�#�7����R�����_��v�����J�,��'5��uH�XB�BIyQ -�zn-�l-A?�Ï���LW$��/�@��?0�n#�l!�ÂC�^��/`�H���	26��Pl��G���"(�8yԿ[�te���]�K��"��ՊnT?{3�����aї��������*;{¨��M���<��������*�PTtʪ�9�%� �ˣy@������X�(�3=T����$%����܋���g����+��-h�7u����:��C���P'	��#��]s�B{����^Zk-�\;���mtq����)�Z{d:U����̞�`49�&vε,�e�\)����[�`�r�uk,�D��yv�a���6�h�5	0��4�ͽ/d|��9jH�?�P/�΢��o�m6��K.-�H"ʖNKťp,�S��`l�/��H�;�*��z�7�%�.D�}G:_���'�`I���=�����M�E�� �'���! !�o�e^ 3�ί	���G�0�$Y?F�$nx�W�J��ZBV�[�yg�c@qT�o)�{O�k%Ƣ�/�i���1�IkH�t����n�$	S�~V��F�ـ�RA��|����笸 �|ۿ�����.��1��Ln|3�!b�|��Ox�
��`�O��S�-"���ʑ�_pSUG�'�`~�+�x܁bN�D6}��_cl��b��k�U6�Nmt:��(cH�&���2#	�I�����2͍|�	*�c�W*��~�3�w�yɘ@G�[RX>���F(g�S��m,�2��e~�m��#(��X4�v�:,F�B@�N�a��П��Y���A��9��{��wW�e�<���2"���n������.g/�א��a�l
����ʹ�qڻ�`)�c�
���}�kɒ2��(�(�Q�����G�y#���$8��ݔo8�I��R+τ��?Ǝ!��
�7i��<��l>�_]^�	 ����F�����t⁻ˤ��?��6<���B�\����;������x�Ꭰ�u6�yYQ*�ѡKs���N>ssD�澐a�U��MCF�4�C�e4��q�1wh�9l�[��D��k�~G�@?U,_�X�`��i� n`��~+9�vƴQ����b{K�Bo_�����[�=����p}7�D^�� ` �?Z�����	��V�h(�񨺅�T���W�gWQ��EPq�l��m[���h��B�j	��Q~� Ł4�Йa�Y#�A{�a'^8Y����STB�6��ɕ���6����:���PgOY���.�\8��ʦ���6h�[����Gd�Y����;���j�~��	 U�ܷ:�G����Z�F��F��4�u|E��t�3�po�nTYf��0��dI�'=(���u��S��nV�;  
���a����3!���D7�2�]J��*�����|It�82D/ӥ�:'�x�Y�)�%�E�&o\5h�䳎�#�j
�������e힭�v�����6W�;�=�\L���(u�mR���0lV�Z�@�i�M����M��~0ۙRb�����
����;[�t�R��?�"��`{� ��(w���������]����}�3� ���;-R�����2�5��\��={��Ҧ҇A��}p��i4�f��Vӱ$��r�/���Q�hk���0�V�c�vR`���%i�/Ëh��V�����b�s��g܁���-y��Ř��g��ׯ�qB�T��v��e�qU��Xܝ�e%� �.������ߘ�O�.8���Î_���8���U�1�H���w��a�ϣ�6�5�d���0ba��S����X���������&����cuJ�(����I�������$�R�W�}Gsd)�r�Rd[9�����vc�Щ���������_=^X���w�7�LP<R�Zm�:��eڊ�ח�k�|y����G��of�|�x	�YD��g��gM(Q�`!�\��.�BI6Պ��+�x�'q;���SI�2O�$�xd���j�#~��װoDk���S�!����ü���EmvFE��ϣ��R�м..;�r�}I�]��)~2q7i14Yr�<��P�������H���Vו�1��u?�%��K��Ac�,���O��R1�0���fZa �t�|�	��Ma��˲4ڄ��0S�^����_�ة��(���:�y�J�Ŭ��;K���ce�2r�P��u('�$����d9�$��ѦX��+)ү�1�g$@ٔ��~46#,v��^�իA�{mi�à�\p�W ooU��6�
-U!f���}3U4������$(d��2\{�>x��$c�˱g3�����;�f��l�!��C�l|=w�;�d��=E�C�j�N�\�u��c�;�*��ê�6�Ç��M�9�mL���C��׮Z����U���T�E�Z�+��v�]_�y�Z�p��8pÎ�-������C�a�e�h����/���t��̼�H�O�O���tz"�("�&͓1����i�C�,�6_N�Q�dw��C�ݞ`�R��,,��
%�a�g���&yJpu�w]p�^�ا�7�Գ�-�Uy?~=�hV ��&d���A���_/�cE	��X2��V:ݠ����.9��x��ن$�E����W�5L]W`�d�xo'��٩��m9JD_�lE�4@�zK
 ����h��㽗��5Iw�ՉJ���8{H����8�l�-�E����tƅ�=V��.��k+[�g�(����9��+W��5I4΂�~�F��)�&��z�����W$��{��vX>��SIMh�3;�)׀���A��ֻ�Z��-�)��,nf�����'�-v���4A�v�y��P�w����V�m �����"ʶ/��G��ا���ڔ?�#]���Ӝjr�#(��d��L4�ldo��E�(�U���#z�?�\݀Q>� �B����"%vT]��씙1����e$N,���)����]��E�ç� �N趢i��vu2�����P��3�k���.��F�8*�>s��^%%�H��nti��8��<�i@�7k��s�� ���*@�J��1�Ҡ��zt��� �D��L?����G�A��֧$]�����W9c�|1����f�&�8璜�G�ή����, LF&�b�$�۸u�5���T{/�1�����b<0�i��X_!pW�o{��>�nXv�K�8��n��^b��m�K���K1E�ټ?U��@'o�t�-!3b�q�O\�LIA��x��������띞�˟5s2:D�gLKY�.����LV�%��4�^���)��t�G  *��.~2B�.��.D��|;cWu����>�������z1�i��$�K����{�|�K�?���#����G�&v��=ӽ�&��&T�-�V|�n�I�wQ���������Gw��D� �?Q�p!�X�-E�w�Ǖ��@�X�ћ1�{���Z8y%� f+�� m��������6;��$kd�?�ax����"���afY}��ک�� �2���s�ww��c�d1���pĈ�l���Lj\���f6b�؁�'���:_u���4�T�K�;��M�T�#V����@��FxT�n�>1eJom���wL|o�Y�y_L!ƗO�1�4���qп)�_�n�`��')R�#}���C� �5c�8HBI�i�c�gb`�~}A<)Glg�.���F����,���蜭����Z_]���o����8���J��i�ˮ&�'~�޴u��o�5F�XJ�ei-� ���q~B��?��]�S%a=����j���!�r��S���{�C�9�"�M+q�Z��\�!�@�EB��Љ���h�E�D^���<�5`�������"'F���6=Ǐ�p|[�<�0�����$k�jg�)����I���L�l�d/������Јcʖ��˄�����NF�Ż����Ml�	�by��,*�)zmi�F�	�"E�z�h�)L���:S�T��X�G�`�y	I�(����`�k�2Q �l�k�i)��)֬��j�V�W�v�PG����!0�rYn+~)z��,E� W�Ȱ&��B`�	��o�x2�!��=;������Q��\�T�ˑ��͞��T��#�F��y�u	]G<�Kq�6B�E��R�^�LA�ۈ�W��*
��X/_X/�� ���a|`��T�,��>�wXX�D7 �%e���������eRգ��h�!��Y�����Y�-9. 2�M�B�EX��VYF�D^���/��jJ���v:Jc�9�����V�ȥt��&�9z�<Ff���Zӫ�T��R�`�[%HTpu���ߨ5�!h��4!}�nF�,����Y�+���!�&\0�y��3�yٖy��b,_�6(��u��#�J㪏�l,��<�	U;���C����|��g��?B
-��{R���R���0?",�,��Mp�Dcx�{��-�$V�;��}��H��-���m�;�T����D,��i�t�����H�L���| "`B�ɩ򀨥�[X�Ȃi�W����5\;}2��
,��pib����lV��P����	��©2��+�����\sT4,���V�M� Lר��A9ATW��ǥ��/k�'�m�)��D��g��l;�dݍ�
�x{\g��^�F<�2�s������7�(������R]��e3=�����߆���*z�m���C�:�tk7a@x��g��+��'`��^K�o���T���l�Aã!�~>*�I�Y�)j�*�JlT~`��p�����ڒ�|�M�U1�D�3��@6��4���X �P*�7R�[�\\���� Zg��?� �!���`��d�6�-����O�M�o	w$�8���AH��k��bu� �D���p0�|e�8r���{����Bz�M���3x#_�Y�	�W�oi1�6g.u]�ȕҊe��B����1��k�w�dd�OZ���0Ng����18�ԁH�Ns�;��e��%�Q�HE��q��sM��"w����u���!{�5A/n��
e��ʟ�"�����������]��9�ئ�����em4�4�s{��|sĽ�o�j}]��?��sc��:_���DbG��r8/�j�t��>Mf�x:;�c/���s'U����N��,�l���TW�#~bz�4Ȕ1�Ǹ���`u�=�a�S���5q45X�W�o8��p\��I�]PD�×jY�����е��~-�N�Y�	C��x��,����&s�Fm͘�J�L�Epx*G���Mq�̏��ɔ����L^'�>wř�պ�u�����H_	�=~�`>҈���`��z����5�״4|E�7PL�D^޽��;���FSʳ��含�&�/��t�8�%\���^�/�>O \X|{LA�$>�0C�k<�B�Z���*�)L�DO@��tA��ֶ�����t2������r�J�#�qc`��5�E�U�J׋�|kjv�G@��Y�����"4�~�C�kyL�3�H���cDd��t��eh�,����Kv��+�Y��!z��S!A�(�O��"���N��.Il����>�%3��W[���P|��=*nb�>��C$� �h�v���&��w\Ma�Fs9e�A��$��Ѡ�>�L{�	�i���f��՟�`He���G��|L.��A�x>�'B&Ж�T�1b�D�:��k���8������[�a���$����M����D��� �LZ�3ך������w�Yp.�$�&
�"�G�׬tW�.J�����9��N��O�:����ߦ�z�9t���3��7S���!��ZO�]ٍDc�D��+�O�_�``��,y.o���ئ� ����ē��2��v��lH��n3�g��\+@D M)'CjL� �پ}-�=��U	�3=�ܚa��d"o���?���F�^�MbZ�}̜������+�xQ�$��HK��N��2

)���D�a4yb�`�ƿ`eP��U�ܰv�ҳ��9s�"�3d�S&�<.+#�N�h�4��G��Et���U�<X �$�A�������1��IG�-��CQQ9"tZ' ��!8bZ�H�*z7���&�	�X=���䍬-��O	:��^����#�4�(VQ��Ff+��I(��vIL�BG�A�=-݂���	F�'*����������fE'��.0������z ��"�lF܈�w|�� k����`��
S��[_Ľ
����-f����,�Vɺ]�s�]�����4�dG�O>m)�n�7�{�i�[�5H�(B��������}`���v�%a==�]���4;��EeI�%�y�TN+wJ(�_�6W2��A��SaV�����8�}�\���,t�<C��uR�3Z��!Tx��k�1��u[�#�љ��7���Ws�@��׉DX=��g�Qk���~�z�}E ��'V�P�T
��"'���e�4�e��4.0m��ī^���G	���Z�
�H�4͂8.�7@�݆�{_kԂ��;+:�i?c�6E�Mg�続�De��) �[���ŕ.���g11��l{��j�xj�b&FM�RU󽷙���q��V��4rR�O�5B.6q��J>+�@�i���H�T�-<;���4�O�#������ڗ#!��-�O,��򳚓�6� ��7U��W��w�y��1o��Sw�V8���{Ώ��2A��)�pS7�����zWĉ���χ?~(Q��+�K]G$�dȷD���b��і���Q�|[$���ez��J�Vq4�kzV�MO��b�!Z�j�~����W2+�.ƽ2�}�#6]��?^�;5sYh��'J� ���b����	�����)��^��+W�`D�xB������E#�(�yr�v�ÝOm�թ��c��x�C.����d"�c�����Qm8E� ��s��6A�0��?�VVʹ�ة�?(*��(F�Y㼠�8͢��'� >�
��Ӎ�ց�A��Gh �`V]��&�2��
U���χ�q��q]�,�6�~���9v|!����ڝV��s��3�x���A]�OS�Y���G��o ��[��+͝z^�ɽ�hq�H ᔻ��3^
珝��~�f�K�ѡ3,�ld�A��� ��~G��r>��3��-����,M�z� ��U����*��̕,�4s/d�R���`�RΕc>��"(��=���>$�����Y���<;�Dl<�V -c ]�,xQ�4XMQ��V����>���頉pe���i/��5����% �B�O���6.r�vɏ"�� P.�@l�/��.V�]o��� (ɦ�7|\C�LZ��L�) �ijG��,|����ʬu-2�0o��ɷ����αߍe��P�8��3 �������ni�i�pX	
���@�_��W@�	~���G���d�H��ؗ�t����=Y!�v\�f5DI���r�WQh&�X�U��� .�魨�>l�,��?�X8E� �V��%�?��
l��"�N�E�,�cˌ�Dٕ�״b�?>ӑJ����|7�S���B� $��./��4�]ƪ"����楱�v �Т?�e��rw��o(,n|���z�GŁ	G��<Q<�#��I��ga��(�Q^��$rä�p2�i����=,���������b����/��C��o�Ө;q�{j��H�a"P��-��}G��Sn��i�YĀ�^��\B�H��h��WտC<� ����d,:�|��в+�D��WӢ	Ɇ��0� ð����9(��=���`J.��ev��4�ǡ+Fʻʤ��5�M_9�T������a�b�_�gaoV��K���sm������'X��J�ٟ�r��u�J�)ϗ�����>�3��6 �����l�5�k%�\�����<zM�n�E>�n%>�S�So���~�Q�����,y���<sS	C�B��@K$�Z� ��"��{���Y�E0	�L��P&�Iva0�i̗VA����2b��1��A.��=[��a������$q-���NZ�5��v�ds���?n	����+-��r����V�]z�#�۱d"�KG��?��z�̰)s�[��T�7l/ ��;�v��h�R�O�5����l1A��"3'/�->!��o֟��1	I��96�y���X�K"��qc�����d�	j(��r�rSХ����D�ۋm�M�c!��ɞiD��fR���i��\z�Tw�*�[��y*�^�ǹ�~�l������U�^�UX�a�9\�@EbE+�z��=_�z�2RN�py*T��J�t���dUMS�w��\C�0Y� -KVO �6$cCN\1d�/;�*�C��k�
)^�f3���O!���EP�k��4���aF����8K� �ׄ�KT�b� ��+���;̾�$�J�GEg���-ǚ��r~�t'Ni�%��ED���J��9�$�]q6J�Cͦp���P��M��q��/�ֹ�Z�ڔ�5�U���'���5�]�՜e���orɌ�8J�q@,��f XY���g^��?����8A}�:\
�B��y�����z����[E�ѿ�.׳������XC�"�5�z0R}g�l:��u���� `�+����Ljs��I�D����m�5�#?�<Չv�V�Ze;kJ�VT�����g��x�~�7۵Z��J����+P�f��l�"#�md/L2�_��hH�Z�8dK�+}a��nIi�2��Dd�형X�!�vO7+���\W*my*�����N�oZt��P�AUE��k����y�02͠����y<z��Ph�rĥ��G: �â 6૮K�_T��G���w���.�ar���������`��|釁B�w�
��)����zw��&����xc@�l��K�����6[q���Q Z��\�;��f0�� '*R,C��V�y2E���c�E=�X��+h�8�	7�!�0�լe��3-���oE�0���������3j�����K���N����5���?��n�@B����"Fӥ���Xp��vJ���&��p����X���WU@=��;���h�|�$��TgD��n��!A��$��4�uZ�3��~��Dn��5��y�%k��.����}�O&t}�\%�"����$r�9��E��;t$̘���R߳_'��?�Z��ua���*����\X)���(�7m��$�����ti�]��Z�Xq�
����ų���>��Ȳ+�����]�7t��I����ج9�$�����x�^S�)�k���Q�B~9w��9��rն;����T��nѱ�ю%j��&nܣ6���'�jvh���$�sF<�B#B��F�¢�o=Ő��-�˹[}�I��W��P���7X�7F��6W��0�*���m�5��p�h.n�$?��:w��Ljd���+&��h�� ��*���'&bH�u)P�C��a��e��B\-�JC 1�O��>��<�1I@2Ӂf X� ���w��³g��j��eI2�K�h����.�kӒ�MBvi,^D���1�)	�%p�<= �d���T�O(�z{�L߶g�Q�������VZ(
�fҞ�lI4�!�=��z��2s��y���!�.�*��'�!�#t���L�*t�3�,}�3kM�^t�ݢ�WI"j�9Zt��xF��`����~e�s�	ך�t>nX���{��H:ehה&�#�~_���K�N��dR�˯�s	�Iy�P;W���a�|C���9�T��.�@�m��Hj�v��`
w��
X{r��6�_��0F�u�6:�9^]m.���ڃ���T�,����8��Tڜm\x1�U�I�T�K-2��7�����=��<"(\W���8�Y"�����@�'!���rn�
`�>o^����jP��W��q� �w� �TZXg��B�f ���P2���YZ�=a�hO�S��Ψ�a�?�L�C�l�ԍ!�Z����=��������.���xw�v8�b�Y�G��M��ɋQ$� ��\��y��;T�s t h����6z ��y	|��u����vnN��ZW	^��v�ϭ��4�iy�� 2:&.�Z�?=\���#�Baj�#?��,������{��2��U�;5�呀x�!��0p�֪�����u�cMR�	�<l�`X"�G��8�)j�QWj[�)���oU�W^�tx��'���`u���ن�oR�3t��b;���>H,�A���W�ƻ�y����~,C�D^�x���ɏ8��3�_����봸�ꒌ��~s�à\	u���*s��+I]�ʑ=�*u[��=��\\�}�]f��vRX�%㻅,S�3|s�#��x��ȡ�z�$�9��#�xߧ�q@��!e�!�d{HDfˠ&~õv�ڡ���e��� <��Z��"_k���]�|�-c���-�������3a����V���-��K١�C׳}���i/$�g�{���������ܕ�q�0K��~ƨ�y!�|��ka������OV�#���	j�'E�e��.�@yÇ_�~ȯ���e9��_hHV�S݂��%��+��e���
�����������7��k�S���w�}�x\�ڠ=|`���xF�U���%"���kf]\��U��ٺ`{;9y��5/7��Zp��L����L�F�Sv�0�ܯ�_��a��9.h�9�#C<��y9Xeg�#���"r��9�tI���/e�Łq���s���@�B�����n�?ѣr.�U�+w}��"�MmA
�G��%�>4;�����\$�vjt��ZQiP-^*��H�$�8�ega^�uͮѤ
���އ�r͈xR��,v�߲n�J�����h'��v�+��5�G��qS`�3b�уf���x�ё���&���#k���I�m���#��Ӯ_#XH/��~��㨤`��*��]��$O�`�j}���ǸOH�dO:/��*��C
�Ob�#iIG�p�j+�.sB�fk�X]�'_����:��G�.�j*�{)wT$l���MCUkI�^��nE잧�20�	N�`�5f�`��l��9z�y��p����������`y�q���.�ܚ��b���h�_�c���XG������_�z	�������������uB�q������CF�6&;uA�}�{4[�C�.	�=W��	d,���/O��	����i�!��쳃�\�b ?�$�ǆ�'Ƣ����n൧(:��\�����X�;2���xAΨ,-��\�.���O��������\�zGi��
�����t�Z{6�n�Bga~�k��S���%��4ka[ɲ̃��5�z�����;��C��I�e4W�ɩ3��b�ɛ��Ku�01>�}�rr�*�k[�Z����@�	Ga��-�c�o�*mW�Q�U��l��Ȳ���A$)�ȕW~+���A+���cU4!�Y��}��K���������.*�t��n�3�R�S��fm���te��ȶ�Y'�?��\��㸰�<���$y�M�y�xM���#L7X y���<� 'Q�Rt�X�4���p��J�X7�@�P��d�L�1j	�)��`,�ʟ�P�ŲR�l�l�
^B}ܕl�9ּ�2�ɦǚ%�A#�@U�V$`Yϧ��r�˺@& s8>�HQҺ̍�R�æn����\�v�y�����}�4c��6��e��]�+(���xJ905
��
.����߆�`k��vz�_���ɧ�i����6�����=$v��N�k�ɔ�ܨ)�M%��$-���ѳ$�ӧ���/E�P/O��w�Z�/:99��/!�;�1ι�q?�wW�+@j��R{j���ua��_)�SP���0��@;�A7��3U ��u���J�52M���u�|%��Oe�T���\� T�MXo:��AP꽕F�𖌊f��^�wmT�.���H왯g
$V�(����I�5��'�g�ب�����I-,��0Z�}�)�MhC!�]
�y���`�sԃ2�'���<?���Ŗ-Ҁ=_�&d���.Ue`�������f��[������s#����i{ ,1:�T�WQb����4iB̢�ʁ��+f䶄*�����-�:%�yU��A��+Yt��DT�Q-'�/A�W��Y��;f�ۢ�Ȳɾ����}�2A�lX��U����?��
��1Y��HE�-��A���'"1��k6��[7��mf���:	���gU�K����t�x�|m��N�����NP=��0�v�ꭵ-;�ȩd;|��̑*�܅2��_a��'\'��8��0�E����Z�Ӵ�!��o�s"6R�fw�7�q����L�6�&�����Kνo�[�g�����A����M|^�D_G��4=�;i��*'T���I���t �Wb�jQ��FlXc��l���N$ʁ�NK�_������z1ަ3v���2��hV���wo]����v|&��"��y�b*vc��^t���dR&%�[&���f�m�d�%n�����K��,9��#��ފ9v
W<��wv}�3:�6aşAj.�(!V������ة����غ|G?{�:��Z-�������X��e��IL\ !n��������̀\/%�� (�Y��_E��o��*�F����]�s�dZS{S��W������"��' ^R��Bc�����S$�Nܴ��r��׆�a��9
 �(�E�	ZgL���+f��J���Y��#ǔ_k�@�H�4T��O�L�G��a���lx�ո�\E�Q���%Y���Q�XN.�]���I��&�g�V�T�D�q��B�#�P�4��lM�M�Qla���X��)�l/�ݲ������(3�0�If6x�W��a�^�����/�䔗d���cE8,���ٕ�ԞZ�f�֍a���SX	Ye�"�q�۫V!ɗiL2�WKYhP�q������7u1�T�1Rϓ�A�>�TnQ�8�iO���;*�a�ٜڊk��'�0];�Q�X+�)�/�|Y���j
[[�ؒ+[�51l'2�_y˔3|�ܿ�?�
��FO��O�
��;�#J��x0��3��{L�dM��~�$�Կ�X��bq�Η��ׂ16d��]�8K�.&٤��_�i�[��}�6jR�	�v=C,0W�P>U�TQ���teM���e^�<�/��2�D��ʈ`�.�"υ�t�]go�v2O��T����a��7h�$�W��@ !���p���as;*%���1'˕:��N�{�۟�{ ��bd
��\�Y��/C���W�#Nh<��W���`Iz��f`�#UA�,�:S��#��t=�ɉ�������A��}B�V����ޙT�{��h���XJ�*��h��x肎���P>�צ�	�i$Bf��%G���RQ�+�Y^�X/��t�窌]���Fpx�S:������
VSh�v!p���>�܉6�x�akcNN���ɽ�^a��x��*Z�[�m���g�op�>A`aڽ��������O+�A6������oz��n_���6z�(�0R�xD���q�S@u<���`�����i)�Cq_����#���6C��3�EOg��/t�)�7D���� $�X���BL��,��w��`�hv���p���?-���q`e��_͘	o��S+5A�N��	$�k�MW:��V��r����C��Sq	�J�x�u8�q�� ��ʭ ��NY�l�cԯɝ��a�[������������@�:�pP5�~���ݎ�S��l��-`j���[�^|L�#~�*�JӮ=$�-Ȕ3�|`M�؊+"V��PZ���>B��C'�0٧�Q���|Q��U�ώs���R�%�'r� 4ut���9f�ɩf!��9��Qwcs1'ppp5˨`t#JU-��%S0��{����D�
�����eO�r�n�]�s|H�xa�+�s�z�E�$�K�v4a�Aٕ�O��ک��N�v׹|@wC3g�n����i^�D����"Iܳ��%'�j��0=w��;\�x��a�����@�W��#�h�1�w0��Љ��$������o��neu������Eޫ�-�w������;Ia��yT�T�\�=Xq^K��b��M����jJc|��z}�E7NC��1�_�:]@^}�ß�f};����}�I��^��Z���+��9��L9k����ߜ�ۿ�|
e d;_��]"���;�1��gX�|"�R�Z��'({v�m�	�LnsX�J3n���gg�a������3����R�KA� /������%�@F�SbYߠ�0/^�1�u�bB���sp�:+�	�TWH��u��A��kH�r�8R�m)�xy�)�u<�p�fLm�Ҳ�k$��k�)�^.v�Cc/Y�������h�V�+�U��"�^r6ٰ2:����橌�@��G��+�p`9=pw!@�K5��o�"k�P�Te:�d��a�m�Q��CE:f�U{&��M��!��x}=�:�d��U�(7�ʿ&�>�~%����?�j��\�4�.��Ԇ����`��%{����2��� eƾ������8��j��,��dk���j��z��5�)����!����$<�A�x�rf@�Ñjl�ZAbhS��{��`).�´�"����C�ES�`�k�J�Lc��� "L>�h�-�k|�C�\�}�:&�Z8^�'�ߨ�s��t�rMŞ!�Ή��%f
�v�Ji+ (fu�F	�O�|0z�F�8ޗs[/���m�Q��Ad7kd1�陠;��;,��2=�fx�\}�_�m/��G_(��82����@%`������Tw|n��R��S�L^��r{q+��/�����S�}�*����lVF�b4?�R��b���"']u�#��9R�
J��ѥ��G��O���j�7��i��w����e&��qG��\)�Q�S��g��۱3#v��$���D��2%�T���8-rh��P�^�O���F�U/���EAn7�9Ľ��^�F/�b���5u{+Z��p�s����M�8��P4w;P��I���[�2La���`�Eɒ��������%���O;�����
�*6�"|9|�B {�9hyg�tC��(XZ<��^���Y�[�:�tUG&4�qH������c�@I[�o��ht�X�3�E��2=�%1bX8�d�r���E=�/���G1fo��6���F5���<;���'��s���Lϛ�v��B)#U�������1c���y��J٢>�W���'�28�2����w�.x�F8q
\���6)�qE8I`JLgO�*�@�锘�(��L�|� �7�������LQM��Oυ����chK�c�;�T���`�YXґ�V� �`�Fd,��+���Ji8Ӷu�	�#>]��i ����̅,cvhYCP6�B��89y��Bc��0\u#:��Om��
�����?�ݵϺ��W�y��nO��]�K�\AX�z �����`�Kw�A �tcpp�;��u<�HF`8�*j�Mŉ��n��+y�<�R�8��WLn$2r�����w��\&}��\��lZ�3�q���}���!T& \�t�p;�P�ZMlK��7���^9ɡ3��q��� �;��u^��]+������V��oNv1m�i�g4zº��U��6��GkR.u�l_�dHb��&o;��T�v"$mD���RӰ	l,�&����D��N�m�ݘ0��u�=���zh5��f�eAp},�_2�;�?¯�Uu��N�wgjl]�CXh���&�����DT��K�8c�BFi`�]ϳrZ�	O�)O6��H�K���g��C�]?r�&O���Q����(,�q!�ό�y���n'v��- ��~`�"bTp<� �?���B1���i�F��;G@�^�f��H���Xe*��U�mk�KaU���D���ǉ��a��x/lp��7�N��P���L+|��}�Gœ�ٔ��}�h
2t�A�$=r���<=�"Cr�RC�=���0��l�f;��-�gX�\/�Sc����ƆuV[��A֫@��'���Rh˹!��ayh?�ꃈ�K#����ߔ�"��k�x���j	q��4a�̕!����oIH��Ċ�w˝ڪ�A�ɌX~�V߼�	�d�T�����jRAhu�+���&�S���3֖�%y��G���� uv�������Q�MYz\P�ZP����	D��Z��p{_��)���%�.K�g@�bK	��`&v�6g!B�h0Ubz�p�/�s�$��W��	�2�O��sE�~��ă>�� -�DT���U�*�1������f�u�u��O\z�FuT��ζm���&Q;$~���w?^I�Ȼ�k��L��A�ħH[�v^�h����'-���T��F�2��"�䒡R�V=j�/�y$�(8�ă{���A*ؓ�7���<�^�̍� ���z�N
�ʈdp�ʁ���N�a#�6F��s�������K�L_�S�é!���A���Tz�$1�G�����~G����B��X�e':��&�E�2� �ou�5	.i��Q��&�In�=k=�P4�kW�D�����U]p��u���;J��@�5�7W��i�ˁ�*o؊�)�k5,gQA�,4Z#�8ab�/��l�m�s�6@/)2/ᲊaSܦ�I��vjEP�0��(�B[��e/�7.t񍆽j�j��o�̉1pf��$|"q~g��p7��I=2�����̨6fCU�U����)��,���� Î�C4̩M	�ϸ��,ǚ�B�S����Љw��ѥ�8�?p���k�:��?pM[�\�;�G}��l#W����5u>",%�>�����Xk�
��_�y�u ��چ�]CoGl䛥��M��}oeͤ����M(���Bo|�P�yj�t��$��wD��:��~	�K�l��'�_$}Z���l&�n����ba)�����B��=��
`��YO�Yx�瓡%M��K�7�#��ޕ����|>oc,Q_��.��7��,��԰Hqc\���)��E��� �+��{d�_3'f���F����gH���F��`>/ё�^a��7�D]]rج�'�A:�� |�}x+��ۡԀ�/
evz.8���I��2q<����Ҷ��}m��s�H��S�-4�ս�L�e��;��C���:�s�G�f^�Ws�7ژ��}�Rx')0���a)���Hp��߼5��X�%�QI��g����ڃF6��IC��v���R�~Ŗ�_Q�{��Xc�{ďl+^)}5�y/�Z����n��+ڋ�y#�����~Oq)�Kv������|����@�V�QSf�H�n|�]��	���\m�W��d��6�^V'~��\|��r�"��63&JCs�>{��4l��^\�4�9ާ�M5�A���x櫷�a���B��mU�+	���*P��߅Ƈc���p{�����Aav��y��*��YaSv�דu.t佫��U�L����g�^$H��(�4����*2 ���x����4��0*����V���Z~q?&��Lz�L�H�s빩Ǥ�,m�S�l�B����NR "�*-K_��F�jJϝ2��[�mC
~�ܒ�Q�����.�[�n�w(G���6���d�Q��ɲ̯��+ꔮ�|����km�e����\\q�X*\c�5$� n����� ��V������Ƨ����eHF��@���N��}��(���X�]�j����J�n���m��Z`@l���|<�G��@�r� �'΋_ks{0T�B�.%i$B�ryb^꾇_��Q8�P�K@_�mϒ$���L^W�gI�A��؏��2�����sR6�m�[���3�R����Ii�݆�[����@��YI�f�ol�����PdY�#�9����$�x	D�a��N\b�&�EmH��� �Vw�صQ��)���>F�1<tf5��o�T�j��;�z���(��Z\��>�~@|�WVM!�ٞg�1�Ҭ(yƪq��#�����7Su$�D���F�vN�������G5DH��f�B�m�,�_x<´����M���(�����������[1���;�&�ne�Ql�s}�@�:�w�X�t� ������E��#��y�ÐC. #�)#��	JHg�77td�'��}�:���G&d**Һ�4J��s�f��j�x��B��Ќ��b�˒���?D�zG��I�U��D���l*�2ܚn�"�'�݁��xU�i
��m,a��ڂ���OR��|	���D�d�b�E"��i�p��~0�K �����Hg5:~׹�ݍng�ٛQ�I	��|�jW.�ɬc�Gn�00�k��#��\JPU�k��JHt��c�8�f9�>z�����P�@�w����ĵy��M U��3L�b0^�f�,Q��5�AO��q���\^.��6��x4L �C^ �:Gն�.=M���.��D�n���I������&JÓW:�W�5@.�M"�V�8+�؃���A- ���D|�����<���d��j  '�K�V��v���]��	oJ ��(��a����%����I�0e {8#�(���*�Ҫh�z���[;C8�T���xU��n.|�4L��E��J������1��֢k �n�D��$�7�,�K��	���X�$����I!2fH�VI�\��+��&�%������p�B}!����u�9�_�݋
�N�V�tM������}T;2IU��������QD_��mƺR�I�j�3'����0�{#�a��X$Ȩ���~�iI��S9����K��.�e>o{<�	�����g�b��e���?��s�]A?C#��J��w6��A�"7���������[$fj��+�C0�r�Zs�9'Z=��9�Z��2/m��$�G���u��'�;xK48]-0As%ז�|��!U������2�֔����V��m�ڥ� !2o�0Q�Ӧ˥d�b�cn��O�5�އ3[��{ϔJ_�y���a�N���+/�ed��pj�+�� ]���:������F�eB�'ۃ'j��'p�-b���	X���]��N�e�j��1�h��O���lD�)z2J	
��stp+��oC��+`O:#���pfN�F�dp9�Sb���1u|�\���)s�%!�m�=���f
S��:v��GH^�
lEg���A�c�*"}`��$���'��,��̍��������4��L,¦P;^�7+�X] :#�	��9%?Bl6��� r�f��鍉��LM��Ʉ�ǧ�����ώ;,��SP�-#p�K�S�g��T��	(��)����=RI���m�	9����	l�=,P�;�v��� �k�T��ӯAKȹ*�^�=s��]��g.�M�ԞdAl�
���S#_�x�o����J�Ӯl��,�z��Uh�>$�)�A�`o��8�ߛ������sJ��U����g�8�HC\>��4Y�zOP�T�=�jɛCƬe��;�ٲB�K�Ο��b�g�q��qK޽�s��֊�9v��|�u2K��'�\��?��P�`�&E�*^�ae{��+I��er֥O���n�F}^:��z���>����B[�>�8���1'ߺx8.4�t�s��n�$�
vk�z�eڀl��W|�7��П7��4�|��=U�+#�rJ��NX/`��.]�{��H�K�T�� UD��v@�%)(%�&wɚ�LSE��g�GG�|�2W~\؈�̾��&�Z��s݋:N���m��C"��9<e��d���Z�^7��0�"c�4�\�>_�:������N.�c�^x�um�|�Ҧ��Gq�����8�í����:u|����<�X�ɗX_Mrg����7�_�X��EW+������ؓ"7�Mnw�e�D{d�����[h\�c�Z�Q��Ԣ����E��ht��/ݜA�ϸC�ڠ��
��;e��Xsm��zZE�A�\��y��; ���UD9�p=��|�J�{9>ӂN�A\��:*��Ki4h3�v�N�M�a)pF�(�F�{�d}5c�Q���gK��S5v�4~1]v��ٟ�q��/����3��tR(� r/����O���fS��4���N���"F������L�է������9l��(we^q�QE�Uc��;[a$U�D4�PČ�_�<*�;82]�2����!.SQ�)T��WR��[ϥ=z*�g@e��k����5^[u�_��M��](7Z}�����Zc]�sAW���1�4$1���؍�Ez�-��Y�"��!� �	sR�}q�[����-_�G��5A$�`"x���=R�������v�,�H�c���c+s��1����)$T�W�ߌ�}4�!8.vY)�7�&f� ����$ǅ5$�BM�ݡ�o�E��X�\�W�������� uxi��&��
��ߜ���d���j��\v׳�%K��b=�[3������>��J�H �7�O,g�
�O�h�3d���qhi��*-����>�d��٫'z�6�����l�^5k����6�v3�r&��wH9��M'sX�=���������A�U��\�ٮY�"2�`�S�f�U�5O����"]��[�>�k($*'�m�o*� �̎�Z�:�|=("16��>���AC<��&���0�L���0&�����,R~ ����mh�'��'�uT�n��Ĉ""`'�K-?�����|$�fof��R�<S�.,�4#�
�	|jvs�yy�Ю�SHb��?�P����V�,�r�����D0���s���E��Ϳ�������5�?�۸��5����o�'�����X71Vw�o����Lh2E8��꒤�
�+i`}}X��Yװ;�>�����h����8l���Ja ��]YuG�0�\6X�}��x��۸�x��U��S:gQh^����l
��& ���oH��H�Z�תA� i~��'��92�P���,q��8�]��/��� �QEw�=���m�R�ʏ>�	Q��.\�b��d��C�R9�3w��Coj�S�2s�^���,Lo��6P���$�wgr����6�����-x4yە�c�])�K����G�5]�C?����3���t��k<qa���:qmX|�ơu�2�;�^꘨;�;s��t� �; �9��`=
�'beG�{��A���&��~�q��iEmcoU>�dXh�q~T6�Q�h��Q�R ���7�AA�_��FG�/�t^��K�?[�HcЩe<�E�G޶���<��4A~
#(+LaS��<� �R�y��E�s�9yR�b,�	����Vq�.S�Gz�ʬ�ٓ l�7�Ԫ+V�6}���t�ͺ���E�[�5���&��1mQA&�Ie���c�x%~5!�8$�f��%=�:��֐߇�W�l�VS1�6�cXt4iT���}IԷZ�'(J����K��D��iƒ~u!	Go��'�B����DŦ\.�W���c�2vUޕ��N���P �w��JÎڥ�l�NCK �Ƶ�����ۃ�� �o���<�j��N_�C�B�Q�����<�Zs\	Qs������/A��P���i�"�\^J ��.��x���F]��F.����~�g���D(a6Dy�C��o:)uCl��!��U_�s�ss��뾂��4��	'e.E�K���y\�+���Ë��z^�tt2�4?��q�~Ї68�+���i�W�`}!j��j/�$��鄜��d�g!��]+�T��3F(9q[�a����u��X?��ŋ�WǢ"͑$q�c��a0�ls�K������k�:����Q�։��	����9P��߯0p�K�MCɭ����0�j�{�E�]�ڭO�u�N�E�"�Qq}23d�a1M
̈�[K��(|�t]��:,�"�,��I��o��/�0کrʄoD�aK؎���v)
3��Daȫ�^P$�T�����3b�6B0�@�_N�QgO�F&o�K2�e_��"��*�bz���١K`xۼ�&U�47�l�H��1�������>sv� ��S�tNѸ�I�i,�hC^�u�P-bl�t5?M���B�M��^	�¤;�1i�M��S�O��?�ErhIaf(7!�kQ��0[Wm�:�6D� PkW��@�e��*�����.��>oL
Bڬ�`)����0���
ሮOT�~˫m�����	5�!�)ڰ+�S����g,_�:.]�sڛ�J6O��e�ghk���z%F�|9���$��{��e�bc����\�Az�tuw����C�xpA�w�<����D��j��ſm� *t��a8�xldQi7�_է-�o"���T��3��.�6���1V���'k��f�T���?����Q��2���\�Bxus}��C�
X�Oݗ�$>p���Y�mF����*�kd��HW.�I'5#�$x0/f��������-+���I�+1�OJr[ryư��	��Le�Bt�C0�q`�a 4S�;n��]�8by�n�sWA±�%wa���}V$�ᒯ�{�'��8���β�0Bp�?ò��a�e�*�X>��EƱٍ�ԯ��v$vn��'̎t�q��.�Ze)q3�:���*cZ�>�~�~�e�O�(�gZ�r�!����K��Q]�9��Ah���;B�[�f��U�Y2TC��}:�2u�AN�s�
?H|��O�3�?X�`JT^���߯�' .*|����2���R�,�~���jTQ	�P[L��kؙ�TĬ.q&���#<��~YV�X���h7B�.]m�W���2��X¬|�����M&pt+�ϐo���{�s�=�~�ƈ�9�D��ta� �#��0J'�"��S�մ~u�{��� �g�p�qݖ�je^�K�^�8�Vϟ��Y��n���4�g���+��������G�r�	�r}:vi)^��7��XF�1���D�	�"�IP�=�Қg͉��-���t7�����f�P5�Lz�;���w��\Tc�S{�~6�t��J6�t�ʅ�����ysB�$�k�F|+��������^���$C���T^�l�Vy1�ONiy��%�%�Cg�B��� b�0�vkyyY@��seUJ��������+o92�a�_		��ծ溊�e� �o�C��ƪ!�Q�ff��T]�C�=��,��{/�f���؀�y�&��<.�꿳�{��Ϯ����O��ˁ%ޖ�_DH�.J fM�"�v���9��߻��P.�/-�s��sNmS~�wzx�XWo�9ّJY��e�K�hjY���B����7�&W�Չ�N�Q�I�4�ˠ瀹�+��ɹ"/0;���EW/�(J���jS.8߆r���;��,ڣ��AbM�&�s8�*�IO��̗�l���{��4�*qs��r��ِe�������|]��c�l\�Ss��fS�/�\��1��Z��c�Ѻ����_K`��ɑ������o��dYU7�I�ը�=��N8�`T��c6�œ,`���aAy��wd�#�JK��:X&������. 	��H3�.�����ੈ�Q�KG�p�O&�����+}M�ǩtou�CF�z+{v �R>=p�ӧS�i-���J]0S��4�R`G^	M��A�p��f���s��h�r����*��.䯏��t�����*���V��DE�W�z($��rXpL�z��*��E�'�R�|�uvV-����vuSt�7�/%��������O������8��V��_�OGO���2<~�2$�CQ��2���a�V��M+9־�G��ۃ�HH�H�"|���1�89�o����R�'�?$5�S*����+�#��Ϭ�M�nJ�f)��ٽ�$z�qE�Z�R��3A�:����onvl?$, 0��'��T��)U������m�4��rB�����Z^:3��8K�������~��Xh�$�v�
�PԆ�.ڈ���&1e<=��K��	3bI�ð�����UDB�����wL%(RC$�����#-�2�8�&Ay՛��6G����bKT����h�>��.�G��Yt<�i�s���i�2 �ps�Q8���ԩv��>u&��(�2�W,�.�?b eߙ���3R�O\/���(L�x�W��ѩQB�jj��Z�tD�4�����7b.Yh1<��8L�]�o �l�D��\�>~�s����c���0��7u�=���t��δT������K ���X��y�JF��/�6����D�����O:#�#�Y�*�K��F6����=~D�؉���'hL���#_����jʸ�h X�XG@<��������q����A�=c��'�^�*���6yz��DF�/�×7s���W���(��C�a~��;�̖��s����G���Ҥ@M����`��:L��(��T��P�Q�v���Ig���]����ah�l��;{�F�Jx���5=;G��ՠ�CO(
�Ԣ�X$$�!��v��hK�ٔF��k�ﶘ�WY���D�A�̎V��ymM���<ʧ�{��8W���*�R�i�c��?vr��$6;�������O�.f�Qi������/��Fs=��	�Hp����G]�%��!-gy�,4�VjH��w����R�c%	Y�b|	�%f��^!o*��H��P��i*�H�w�-Gf��6��icd	��>��m�0]@hj*ĝ	i����9$�Y�Z�!J4;z`�*T��/���	;ᓳ.Y'L�+��V��%�=���-�O���A�J�6?����;� �ĸ [Y|��3���P�=�u�g�GێZ���J?��,�~a6�? Ļ���1���6�|B�	�;�3.���]Kb>f�F �&�k�{�
�g}�_1�G��&�P��|��~��Ix9)@~u �9�q����Q��iӓ��#0��� w�C$)�����-�I�v�����)�S�"Q�ې��v��Rպ�V���T��1o�o$�-�ҭ{V��k�PMخ@MAY_��1b )�_��w}x�P4[asd4��1o;����V�o ��@p��u�i���?��s�a0��u���,�;��Re/�j?3wF�`n�o��lQG>J�%��޽ͅ�-���)�8� ��Y�b_�ؖ������F��i�C�tG�"K��̹i!�]�8�E�(;�8Ֆ��0%�옗@�- ��o�ZLH�Avܣ�>�2���s���97��[�_Of�\35�zS�VB�� eJ�).T�95&�:��hpWTM���e7�?̆c��ɯ��m�⿭����b�S���*,�ICr�S���9���ʚd���l��e��<enAč $�iCIi��N�i��eF[ؙr�L�����A���  �@��'"��9%��yM�kIM�J���v�~�2�M��73���t����q�������;�c�
abp���!�!P����m��B�N��M�bDF6,���H˲g�K�Zy��b�Q�عa�e�-�)��Gvd<�i�(dH���֏[ڣ�\���وr���P�%Ϗ�ga�g�=��g+��4y+�H�w�R�_F�S��;��(G��Ո6ݔ�l3�c	�!"�[)`�i����M4��*��C�5��}��*vb(��_��Aj�i1"f��>_�DQ�w3�l����n+=_Ҫ��a�h�;�D]o�~�P[ھ�Q�1�!a�	����o���4�����j�}O��ޅ�;!��(-"T��09��X]X���hY�g> �u+FNۺs��+<��=A^�F8�&�Ep�ˬ�v�1��_ lۊ#��k>z����-�2=0�/wI�S>ICA����2�"����Ŷ��d��Ė��1�S��S���3�YW5Mgg�n�X�>�..�/DĐ��Y)W�ڠ����Y�6Zda��U4�
�ʹ^���ٚ$�����2�tц&G�Pp�~2���N���I���^��[�R5���BOH�(��[��s��k1��n�0SSj+�ff���wԅ�cU�1�_���h}�LXŇ�Jꀨө�Š��4$<���gtO]��N��n�n��sz璲#Ҋ�lo��,�&[)�b3���:�gD��]�~��\� ��BB֔�b.�_K�F?��nHY���rc���T�3��C߭n���� S��"ta;���]W�JЙzd����u�t#H�Oρ�91!1A�VN���S���{\���=�!י�-�5��c����8�Ͻ&�efAg?�7�ʶ���s�Z(K�L�S��M�p���7�pѐ���t����];o�;�����)�y9z�x�"�sx�%i׭�C����o��g�����t>�G����߇�WCξ0.>����."����*x���6�����V2bk��r�H,E������O�M�v�e�]7�T���FK�� T25k7�`��Ig�gg���\�b!5U�m�߿/��V�so̹�P���y������ >��x-j�ZRYNPR�h��A��� -�'D8Q�zV8
0��X�M��q~�BWF�4�F�/d8�N�b�iY�q�� :r����kk0>Ķ����5�v�-��'8f\ E���d}B��8"+]�om�s)u��{q�f,�nA �xc"���<��"X�N�-��ŵ�wBYĶˍ�:x'�On^����v�d3V���9�C���cE|ߕ�I�-�@a����b�jt@�L+t�$|��v?��r��*v����E�u+�&�}�3�D>{��jFb"�/��7�C��L��gph��K̍\�P��$
�&gu q��6W�ڴj���XM��Ty�y�O��� ��DqRQUo���� M�5��ZE�l���yE3u+=���)a���q����r���N�0IR2-����No��0�C�6�x��L�&��hn�]��
����n킂6��YA���	ZT-n>���Wڂk
I�o�r������!1g�o-�R!����&�qf���\ʑ	&�Q�+e���?�"Ʊ���wCᕩ.!j�U�w�;��%����h�6���;2����:��- LlP�����{�X��[+��c��y"�-{s��d�C��s�M�|��n���zZ�k)���^�.�07t�N���+�ǍM��]o|o~!��M�@�sHv�4Y�ۨ7_���h:�1�8|:�Rp���D~Ș�F���pi�e��m^��ȫ 5[a(�*�?[��Q��cZ�SH>��F�����n-�@^s;��f��Y��������	n�w���?�r�V�Sʖ��baѻ.�Zc���+����� Aח[�<��I� �@�s��P��< 
��?�-,S2V(g�;��3��e'W���Y ��آL�T��_���^���
D�:�^�WOĪ��*�_�- i�=�@��� ���X��t�%�ֆ'S}�*}ǆ���X:J�A6�s7���.�&�MԾn�ٹ&]�?z(��ԁ�4X`���#��8�<�N/���4х�#㉌��y������wSk݃�mpi���Բ�gg���0	��7O�v����p'�>gZU�HV�U�y�МhI��R�k�g��$��6bƣ��^�7�O��̕m�ګw<�jeA}�3A��K�7��Ҕf�#�Z�E���bKXè���:���Ϭ��mo����fL8"��R�>���k戣�I�2K�q�P���N��>�1�"�	d؁�m5�0�Q���;N	�!Inb��xA���\\��[������#�`��W3uzp�m"Зf�����C�)�'�5:��'����M�T�bl!�*���7�XGWM�p��
|0�~;1}o^�q��R�D���Je]�zH�ؠwѤJ*6� ���Xޚ!�M��{˪�Dd���35�\Jb�]*���-V�s��&aIJ65twr��v%�՜�#~'E0�MѠ�2��p(f�F"=��!R-�V�HƋ��P�^������C��s��SL�r��7OU����<�����v(���Z���=�ဎ�p�
���CZ��o>�Ιס�����B�aV禮œ��<˴	0Rhb�JW��<����v��=�pzX2g��!Ѽ;+%8�ET���Mb��%��<�H�@�=)���‭������	�d�ܒYl�J��=��*H�y� �u/�.�.�������8���PdoC�qR��p"�`y����~�V:7g1�	W���|M���v�%/Nĳ�i�Ы��kT��wr<�N[Ǩ��+m�:��7�{H슻l|w�p$���9ݕQL��5jݎ�7�`˷�iP`�]��H�3Q��;�",3�&N[Ki.]"�!=l����=�qsi�s'��QQ�u��n�̟n��6K�M�-[Igkr^�K1Ƀt�D�3���B��B��)�j����[N�^1xO�C��/�M�-�A����L=���bo��'ףإl6� ��t\�0}WƟ8�C��hm��
#���
G��ܜ�N�G��u�|�-LZtA�gq����Kץ���a'}I�v����m|�z+��j��E	�vU[I�V���nc Ĥ�9�b��O�1;��E�K??%0��,h�~8zH~�O#�?�W)>𴐛��t������Ke�$ɝ���ܵ�ƩD��c�[^ �r�bHc��K�[�<���=��КgL�:6ɨ.
��!�݊�.� �\�,�_��s`�x���3�Q�.ئG��Q�;���N����w�X�ݿ�[;x�~�:HG8��!�:UC���0&S}�)v�����)�#�`��?C�XyN��Hl{;�ɷ���)��t�Ќ�G�G�����:XQk?>�i}��v��`�R;��Nq���e[��<�M�n@�mY+z��~%�4��ˁ<��P�TLy�ij���N{�9�p����C�����f	G+z�B'	�@Ly�Җ�=�t��Aŀ�F�T����>��B~'^H�ܣ�B��1���Z��:ɳ6��b�:Cv�\ŚwEN`�L�c�ea7_a��
�Q�8���DH8W�uӒ���.ޱ
Li����AvJ�ʸ��� �Y���f����2'JX���9��CQ#P�o,��M��q���5��=4+��I�X���k��:���a��*�-}�]�:`���
o�`x��\��C���i�s>3W�\�ĕx�R��9NN췋��z�)Kǂp��d��O>�pl����
�V/�y��,K�z�E*;�$�c���[+ ��{]�c�B���X����Tu���;�3!c���=�y�T��E�!ngˈ����W,��eB��<�Wc#d�8r�Tng46Iĉt��u�2���ͷ�@���ұ�R�j�<�σl��DS��`eU�,����g���G����ڧ�jO�ʍu��K���BT2&���};���%���a�}�\�Ab?<*��R�S��hV!Grx�!EՔ���4S�P��GY(U�s$;}�Ea�3g꓍qj1�p���>�2!AZ
J����0 у�9e{�;�����w
2#	r(Oia�5v���H2h����g�6��Q��O���T�ͯf�܁���%
3(��
Y���冒d�{E�cH��h���g��ғ>$�&��2�w���4�N�4�4Gb��T�1/����ۮ,��b�H�  ��|�N����e�$'�a���ᐾ��mC��7��ٳxK�S55D�NlB�ӛӖ��
��`h��b���}Y��%�xqM;P�����W�#���ʅ ���������1��B<�-�疙��s�J����E�=����;md��q����K2���Ӌ#1Ц�*`���O���9�.	�IU��������o� ��cٜ��mK�0��AZЪһP{����-,�lfAzf�\U3��T�g�u�R��m��!�c�4W����C��� ��V�/��zC�-O?t۹�hqpM��{3�Su�N����KF��yu��m$��+\i�bK� ��a��U:o���_���^Oyg�裻��n��>@#�O�"Eê��b0�6����F�	���
�+��}6��|�zDa�QK�$l�*�u;�}�{(�,���F����+���ta��R��;�ݥgMi���'վ����*�{��nVg�v�c�#H�>9I�|-��H~��\�8%
^�9���YS0!����M����i�J���x���> s���(1���@��p�d6�A�B���)��9͵G�J;F��R	L��N<�Q:�\�L�*D�?�p�H+s�m�XZw%\��{O�i�;Y|�����s6����_������]�d5�������t���NF2��� ��6 �sŭ����D�u�b��ۓ��X�6�D�Ss���Z��r��V���k@벨1��h�9�� ���zSκ�����L��8���1���&�h�<�g��ц�E�}1<�hNvi�l������'
�Nc���3T���3��Y���\	y��ȍa�`w��O�*<���z�JxQ-[*/���X�^��Ye�N����5F@t�C�Ar<��?	tTXo<C�wW��	~�i0^]1/�o9�@Bgϣ����6ŵf��括J5s1^̾�"���8�b[=���
s0H��I�a�5X�$hO8Ee8|ޏ+���$z���C�=jx�h������x�|V�	��a�7������b88H]�&��!S��V�Z.<6*^��zY�ϲ�+IU�K�GE��qh���ԧ�Ɩzڥ_�(N��UqW�����r�;ɿ�%ZU���4�6z��i�Ӝ���k�<��VN=P.}W�"naW�F$e	X~N7�υ�����Db���T}4�o�����+}M�W��F<�y	��3��~c�@D5vc���JJ5�P�hƝ"�j?8_wZ���ӫ�C�бz��e����
qx�S�ҥ��O=K`}�ң����.�3� �Rn;t}b�fy�&�h6)�[��\I�z��F���	sJ�2'Ͷ��նAyO2[�͈:��cS$��Ym4%����A���~ćwP�e3���mB"�`I�v�0���$+�b�֭SlZh��t�ڪ��iO`
��*{��������A����Lf�7A8���4���?��b�D*x�i{�p �C�BP�ۄS�N�4�oS��Ci���ۻfc�-%&T�d�Ek!K8H���)��ň���=!}�@�����%���;N2&��<�"B�o���	Y��&�;�t%����{N�a����,T��K�7 ���W;UA	����oZ\��q~����_~+�V�1<뙎�m�I��CӄPi��~���m;h��hN^[����$	�Ē�|)�9���w��gʘ;�� �����R�����%M���=���t6	Zdr�x���`(�y�(Y��p�0�r�� ����dF��V��a����dhN-����L�t�e؋w��D#���z�|D$�:���_��|D	�iCS���As2��F[.�C�����T�_��p݂�:�CyU��C���07�` t�j�H���Š,dC �(�� #��?�"��6+�+6��A	eP+���?G�(��{�+�r/Ȣ/��ɠ5K����B��j��K��P[�K-���?��#�%��AFLY9=�=��ѷq
�u[�ѭؾ� ��cm���@��e}I�Aէ���2�X߻;��ρ�ܨ���ޅ1M�gy�����5���!r&@1/�-$p@.5���P^�i�~M׺+�k��"� ~�~����13.�g�N�O�+x��׸3�m
���B���瀶���������Z���C��Y�T=��.B���_Վ�~ym\�u*]�ʥ;֣�Z�&e�����ht�˾'~Kt\�N#�kL��Qf�	S؅ւq��Wky���s�[6���p��F!,ʿ��\�����I�����m�J��/�qU/H�G�*�[��EuSɩՕU����x�(0�0�[ޚ�˃Q�4�"?�Գn��^�G�2=Dr,u�R��]�Z�}�Sj��h�{P�S��ԕ���g8}�=�b*SMvI~S�ݻH����4�(3�r�X���eh���-G�$�LO��[�q����>ڳ�g	0㷣��',����>r���5��F�8~�|��<��W1E@��D�BG�ѻ8=��}|#�l�P@�nY�� ��*�~�݄,�8f&�ִ��ܮ���?��JO ��ーK�H���@!1�E6�9:J�="s�}D�!�|�ik� 7���1O��]�8;U���'�i�V6��(��
��(����.�E܋����ѯ,�:8.co��_���"/����)=I��4g#��Qi����{�����d)���W����th��VT�O]�&���2b��)��ѡ��!?���������h��u�&�a��Y���J4�1���?\-D��5Ց���jk����q�P+��b��=�Ο�+��� ���J���p~lP��(�Sȝ�n	kO���Z�?��Jb�Jʅ��Hw�K�d�ͳ��ź��2~��(^Y�������tt�GL3r�T�c����b�	����Z���ˋ<��^޵�nɂP������^�q�����?[CbW�H�J
�����@e���@�O�F� �Q�b��}ۄ��p!H��F�.�wrQ>1�bO���V'$:񷰊�j]�s8�f�ɂ�U�K�������}ܻP�qV�s���n��x�࿬Q�	2�F�t��u�\�K.���Kv�]ǝ����me���~ÛLk�Q�0z�`̲4�����&���0�iζ�)~�v��c� ��+�,�&�(_
=�%V-�T}󹍀��[��KK\�����gYq�A,L�&��ɯ� �n[�2�:XQ��EI���\;߇_(B���x������¼�i���=ȯ#��.�t�q5�T	���Ē�X����UB :3�gJ���� �5��g~�`Q`�����7�n0)�`��YI��Ś�x`�N�B��44۔R��z-���'�k�51�=��t��oJj�%�2���&���ˊ���fzZطpEL��S�.�<
Y8�'��Ε�}��U�y�֓������&%��_�(-�-@=N�{C�#�(s��g�y��,�����=N��=4%��p0�i���픐��}Ó)��KX�^<����V1%�g;8���U��7�,&��nц�h��My}E��MN�R\H�Y�g_]ւ�^���;,=��X��/Jl9rK~�|В��yE1[6Y(DɪŪ��,.w�TH&-���Z�X��DA��2�8��JE�z.5T��bRl�uQ@����ñͬ���)�8�/��z�b��ڀ R���F����c�1c咐r�lP��L�Լ��F[1����՟
�� �v����>z1cX:i��@cZ\��6
Qe2���� �¨���Ȱq�H��h5OrHB+I	�vj,�����
u��ݠ�W���PzX�}�py�j�)H��#�R��_�}p@톯��c��G�ɀ�H#�����_�0�3aUg��p���tƐ��N�5�bGX�������z��1a20I��/&��F�M�A�#�D���0e�yi�Պ��w�MӚĸX�VJ��<�^��*?w��I.D�q�xt&6+�֖��X�U���4)/�����m�n �d��y!��a�P4�F�`d�.�ڥ�tB��^���[=�����ݞ�Sx,
|Um�0�2õ���c3p�����FtiAN��Y�skj{�L|���(��u���`v߈"g@i�&B�?�H� �y0.��C8��	\=�}3!K�/�!�+P;�h�6�]��1b�p�@"Y�ޔ�6S��w{�y����lp��aY�n9����[�@
B�����<�C)��v���N:��z�

�}u\��9�W�K�ܾɩ����$hYSV�ۄ?�A՝|�k�DK�U��;s���|r<^N�~U�o(����[Ҿ6�Ǌ2�?��bI�؍�w_�������$)��]��d>�y��b�]��`�.�* �Y�����U-�u��A܇ɧܼ\�{��wW�q+���q䴘lmjU%s�X�C�r]��,u�!�_��h��.�i`��l!�:hSd,����e1`�J���n,��ΌM�"^�1�&��7u�1���KE�������W�M����4��1�~�|�����*d�6�·Br����KY)f];��Ƃ���U��t�DK�s� �И=�ؼǿP�:a�I
΍��NM�+�H��7{e%L*SN�0�DQjL:G��hU/	���W�`���x y	dN��2E�13͙�D-�����s����څ�S�������}0�&b�8���~���fT8��Q\�_.)՛��|�NgO��|��@�l�?l#>7`�q��=Z�?(&Pb�I�^q�=m��gD �j�ϧ��+/ᎎ �b���?�C�׿��C�*Х?N�E���5�~�T4�װ��~ȓ��=��i��x������K��K0XںI�val��Kh	;g���^�&�q7.�/�G(p������擄�Gc�.5��^P�8� �=mP�u�-�����Y���_L��	z9��Kq2
�Ta�M#� Xi��3���@��2�(�g����Ν4���2D	E��@�̦d�%���o*�2��5ϫ�fС��WTp�A'���G�k8�1j�Ǵ5Gf�s��8{1F"�*����~t����$5�nbG˴�x����,������1>�L��dS��C���"NB����-Lyv~#ݥbH���a��!��s&�����O
?����O��[ѹ�@CE]|8�2P_�C����E�M��`%��h��P�(Z��N���v`��,�5@X8zLw��)'�m �oA��?g@򠥉����A�V��}�.� 5���q���&�K�z
�@�������iҨ��9L#;�/o`ܜ�y�� %��e�w���&��hdQ~Vns\e��G��O5��Hn�ZFi�DC�f�k{ Q
�)�Z��2}`�m!���F;	0���h�<��AY�]X�@�ͫgM��Rk��eo�S�{/�Q��;��Y2���9�P��:�7����nv��:���r��~�-�;y-LhIi�NfE�Uh�����G�zs&ܢƍ횹�O��Q���@ܱ^2b�fq_��'x���n�v�TC]@�����a�˚��9��8�hKA�O���-6���Ԫ <`8��{��h�"���܄n���ꮯc�>0-4C��&g��D���\�Q,1��P
�c�n�����gCn��]��f� �ǹ���	�0�v��Db����'}\ɫ����AZ�P|*��;o�_��20ΌD�*[��bm�&=J��0B�,�	��,�����yUn�_� f��6ea���z����<sR.o�",�zԧ�����='3!�r�p��z���u�����Ȭ�|>��M�ٺ9c{���@�)NVXvM�_�#f�Fz�xd�:�5�16���!�#h�~��/��08Ԕ"X:��}���V��gH�ꂜLf01
".�:��c�J���9�x+��e�I2��&�yb�Q;�=I�8�i�v�,�d�hGg��W�$B �x���ѷ6U,�,����h�P쾜�� �AsNO�!���b�x�BN��bK�%�:��I�;�����:��* }�ğ�e��,ZX_��OJ�?��`{��T�u�:��*&�K�E2�v3m���Xvk[2;����J0��=>����l8�y����y���R��~'��+���"j�:Ϊ�7�K�䉨��v��;��J~B�]�|N�Z۷�)�.�ɧ�%x�v�O��ֳ��wFr�O{����&1��>��^�q�]qx�2�
#׸%���Y����A���Wġ5�����$�LJ���x���푉 �w��%�Z���V%������p��)�R�1�̰_H�����T�Q�]r��_�v�ۃ������j����6/'�#�=������zj�6��ɛj��w�i��ai�x��� �'K�H����D�00��V8���D�\`z<�;�(0�	e`�p/�Awl����
r���J���87)����K����,��=�/��!��]68j`�IʁͶ�H|n@���'�r��l�P�hP']{P'�R�[�%����hj�oM��jv��b��ai�������(,���
��'M�r�i�|�iŢ�A��H�׼+�:�YqeF|њ�}���
?�����mi�μ:EvG�. B��L"{�E�Q�;z������wz�nO��-L�<���z� ������J�`�KQ
�k"E�-�=Ϯj 6��L8^�.q�����ޟv]����ı'&9t�ST��f?yA��`X%�h�t*+��O^a���3���1$.`|J`z@�B;d����M�g��
�S��%WlҊWuH�*<5��-�����!�(����|�%���c �%�@g��.F�K2�`(���t��јD�e"POH�ύ�zY������7ͷ!��9��q[E����,k� "�����Y��T6/t*�"��ꉂ@KQRY��:65�M�
�Wx\���c�G�ك� ��:6��_l�r�VV��+%n��M�����Jh�=[	˦����띠�s<M��P�淇d�:�騐���%1fN�5���A�$�Ch��(+F�e7��z�Dz�QO�<�7��Gf}MW�k���x��Dр��6�ǌ����hSU�iȪЛ��\@1���4�;�
�$^�]%-������v�������7�dF��-4u�C��22;���g(7!.4Zs
���T�O�8ĸfǱ(C�b�pO���ȡJ||u�o����A,}u|�MR��/!�,��\3`�܋_����Ѫ��C�&2w�:�l�3\Kj�C�a���cK�z�~y��\�ݭ#�dhS��+z������?�+yT�}ނLB�w��^�tf"U[%�Ջ�+X�01�ߗY�l���A�W�k����O�HDKxy�kHB�N���~���N�ӄ��!>
e�0���M7��
~��?	��u�]���d���|E��O+�C$%v�M���Ͼ�K��%�J3�j�z�V1�ߓ�P 
J3`�+�5�J�l;f:�%��Fٮ�ʣ����y0eQF��;}c�S��,�p����x�X�^5N��x��l>,�𕽢^Xz�#&�߻D0���Ϥ�s� �s�P� J�K:%�Ťrʁd�G���+�-���W?J��r/]�� ��Ãt�P��.��Ě�O5�@��S����pE�~��T]�NFT��#'�X̋vtO*�`�,�e-Z�0�cr��8���)�oW������7��T���=�c"��b!2���t��S9�O3� ����림�A^�Q��
g$4�j��p�F��p+�[�a�	2@��ARS�r烙���[�\z�e��,�'��;g��u�ɥE��>�t��f0���	R<�d�J�++�XR���Ag�tI�D�c'2�?�N��z̋�{���5j�o�#n)��j��;��G9�|�5I�BI(�h W����9L/�ND�ܱ��h�����qbY>�H�[��>B=���Gװ� �}8��D޾���'�$��m%4~SeT��)��%G�/�tubMb:i�=�߹� ��=����� ��Y�F|�m�a�����p���#�e�Kj^J��U��o'/�mb��OA���<�gɸmk����78������ ��F;���*����ֻ�<Ȧ��{�����E3؟���Mq�P��6-�qu�zH���?'0e�Y����P��B�&>�ݩ��5�.9n�G��MfH���U�ag3��bXТ�y�!Y��ۅ��Jm͟����_�f� �O�O��ZO�i�����,r�:�A���^�˕��Wi�*�-(��/e�4M�M��� �bx��@B���G/5@K����� �s=��6f]5��m���i�\�ӹ����ƞ�(e��!������@kkn89R���A�KZ��P��؝��.A��n" �<�xO�J�MJ��9�w<Z�	^�O�x~G� B�gg�{������	��$�O����|Ł��tԚ$e�������{`����a�'�p��o��=2s;�E����b�(���^�Lx�{{�BYX�����푸ZO������_u,Laj�?��|�W�V̱��F��r�H�����J��>d��OY
Av�bl��#Ts+��Z�KE#�8�jY�
�^����j����h��C&W4�>�<0/��ѵ�ߢ+��i�_l�$bU50�[ǲ�������EI��?c�:�:&aߺ�p�Sk{�����ǈ�h;���D�C]6�֣���)0���o��'���˒Z#���)��	�.d�rδ�1#Mhtm�D����b���e&=Nm��B
�f�p�u�O��д'�yK��*���)[�%2%f�������g,D_��N7�����};a�=�8���&���.$ib���Ͳ����}��U�����؟(��x��},U���1g��eݟ&|��R��B�F��0T��+��|����J��c�nsO��F�JZ� ���@f٧�>��(�������K�H���{|sÑ��>x�Ze�H��X��ky7w�q�is}*���'���v�C;�U�G�A��L���M�G�.���Qa��6^xH�h]�P�h�S��i��-+z��bK�a���U ��ǈ\݈$|Xq�%,9���+:m��pL�Ax�<*m���uIV%=O�a�6���x�da�㗣 �x�ΰr@��(l%�'�]AO���,
ͺH;V>����b@����iA�8֙_��K[J�Njc�����!Ԛs�XſT�������h�21Ui����GT>�B����wd��QAh��u7j��u�p_4*�99;�㢧�m��a��19;a�!}��J%��p�����᯦ΘH������XҼ��'ԬH O-iV�D<ɤUI<����M'�aV��&P&�i�{�<^�k=��C����d��>�f�!���S>Jr��^��~!�lT�.1����&/�l�O��d:@�^)��40Div߉1b�Dyhyo�NGL2i��(�ʹ��$�z�6 ��ޅt:|st{�'���|Z� �n���V[���Q^T[�cGo�v�%&�:�p�Ϣ��\	���n����k!����a��$*{M3�����J�#�c
���q�b��Inug�I�&��_��ҌT,��ߥ5��/,��eq����Ix���b����K�@������Z��:�?��2���sJ�]Կ��Y>v���)ꡲ�hN���h�xMC����z�������!���w�"�~�L!n�̻����a�x�%�Bm�3H&��d�gN{6z��\�N���� `��X�[����q�	� ��T}F |9��1���\ lyX��tB��p8�sX��U� P�@��72;��. a�k|f�N��cL�q��ܕO��I}O��a�Q+u! ��(~3>NTNbz�X����L"��V&���.xm�\����r����{���àZ��:��<�Nu9�_�����k�p'���[2`_$�W29=�+��9���^v��u����j��,�"'��|&���az���0��G̛[���m6-�����6TU�v�s�_�٢�6o�u�.1VB?�5��s��-{��.o�ַ)���9�V 	���Y`w�F
�$.x�9C����Tz��+;�H��U���Z��6QKq�O{���Ly(��VQ"Л���Ƭ4~ê�m�z�YQ}JX  �Ѯ0=#]�2z�d���i��4��<�<q�%+�
�GŁ�1̗U��|��v{�D�����(4��Ƶ��k�G���0���CrNY*��V�n%�pX_R�VMH<)��@�[Џo��I�� as [E{@��X���nw/|.��4r|7����>Bɼ�-�m��kR�f��c�K��O���_��}5 "�_o����뀟&e�c��䠽��J����4o��If�Q�ŉj�����,l�q_ʷ�|5�S��E�_8D���#D��G���	y��Bqz3�_��n��~OVk7C��� �kN|W����#4�.)�\4�/X�}?�	
��®{�>R�T"~�e��X|�(i���u�ٟ$�$oᄧ��֨�WN�@�l7��r��aӍ�&h�����6���#��OG����颙2S�"Q�����`��b�O�X�d�y�3�؋��4"���a�=���ͬ�I>�ɭ��� Ψ g58�B��:���/g��q:�'Qn��";�4�r�)��T�E�+��R�.�&��#1���g7:/r���`�J}qn(��"je��ko]�\a+d��H���C!7�ܑ���#TE�E��YH?��V�����5���>��[���0�7؏�T:���zg7��K��!GzoDo�k�s�&��#:���$��)$̓��*IA}4��z�%�z;�8��7�՗����_Q��~/ɩ@�,а~���=�Z ��)6 �\y�K��Y@Ho�����fI���&�z�ߩ<Ol6�Qx��u��VqXPW�%�u��l��b�≏v �=���^'r�ڝ�l\����F1I,"XӹyC��HZ��A��dR�ᑾH���55L�l��DF����g�ql�Թ����ϝ�QQ��rl.��ݐ��,��t�Zb.}��*w��	�q�5`����'��8�LvgGr`.*�J5A]� �7ɞ�T�bߘQ�
U)	�����-B@3�¿�䘏����ƶ���֑�>�[�|[����� 3��,a�Y5�j��4{@r ��k�c�͇�m>�0�v�%����7GUX�9!A^ �6�*m�~e���@1܊,�mי6�C����ae�TWĖ`ߩ�����,R�^`o��i/��NΪ/�C� ��{h�����퍭H����<ʷ����������#�9�?�6$1��l�>���u�|�c�%a�,�!��E�챋K�
��Ge�!����Oꕖ��y��y<��I˝\��4��jbDw	�by"��/O����y��
K�U*��RX�oz���K(z�	���C=�N���O����� �ݞֳ�#*��O�Y�#>@����\��T�N
�Qc���A~�c&�T��fn;��&?I)�̚Q�lD�N��u�
��qV����/"�S�+����|��t�*3�*��FOj���P~��0���]��Dߦy�,��`>��\ȴ��Gn����֘��4������' ��'9r��מ0|�f��#�'��%�qY�6�h��Y���jc4GA2&�@��	>p�M�`h��d?��B�P�=�?�˺s���*L�8�՗S$����2�D>�$ۂ5O�P ��zn�H��c�^���F�G�|��z�<vw���yʕl2rCơ]9s����h�	�5�B��c�2�߳�͇�U��@|����P�>K�\�ʉ�o�LZH�:��
3�SÊ 9g>��,")YE.���>�d*�k,�m�������c�
ߪ
E�ƿ�)f���S�9x�&�Gs2�q%V���ڿ����o�L�6I�$� ���`�(��_U
5�#�j���~$)�y���Q&GY!ț�c-�X+.�o�6*�)�z�[r�[�]r�n��a�9�z�M�K���J��aI٭;���	���{�6���^��)�2�g�������즖ʯ��]&%K\c���v"o�)�x��n#�P��,�u5!��8m���O>g�M���(&T����P�F��A]�(���گ�{B�<#��n�g@��<�j� ��9�,�?��(r���,���s�B90���� ��@Re�=㽗$���������׺~�>����ǘv��2X�Al�7�A[����h3K�{+c�B�x��KN^��-	�itIT�4J�t��W84je��رPM�0�D�K�D}�{~a�R|��� <}i$��GW�^���o����v��e��pmoNZ�[�!4I.�%��A��B��>��z6�s��c7��R��dZ��|w$r󩰻�c��R}'l~�o����q���;GX��T��[�ӆ���e%�,=��n���-��=�v�r\PI��8���A�e�.�E�"%�P���B",��oz��z��#�}w��7ߢ|��~���a���y�Zsr��S���	���t-n��Z1�����]M����S�6���$g)�Kj{r/��� �an)fȈ��D0���T�+�S�b�X|��a�<>���h�8�7����y�[���v�و�|i3�'�����7�O~gAq�LKX���w��}5J�Z,^�7u��[��}b}nK�[�'8p4n������&)-�8�(���8�S˵�2L���%�2����jn��jz��K7C��$}��7�L ���S(OR�V	p'�V�����Q ��Ϛ�Q��Ű��G��:�H.�_��(��P:� U�E�ڌQۖ�?eu����ķo&��V0��W�tx�S%�Sjn� ���SZ�SrK:�ں���=��(Y��ٷB���x,��1��=F��@�Je��(����E�jR�&�n>mh-�D�\�(.^�|ġ.�8a�׽h�ЍRb� ?�C�������_d�}�~�j��Y�No��
0{ŃXԻ�"��A��ޚo��[M:�}B\��@�'^��csi&)���
o�
��ި	F�-�urD��6�aC�z2��eGI�Z��:Cm4U����N��1��7P��6������X���v)#��Ӏ�3q����^��
���@|}ǝ?L�뱉��O ̆:h�bl{���W��9�uo�����r�,���-ۙZ眡�,��H� ]���
~mp�8ǚ=>}Gi��,KubHJ���9�W�5}"���zA8���T��/�嶡N�ڶ�����G�[������ b�t��H��ı��p����'=S�����Fw�%l��\i�� ��6"X�{���ˇͰ�ݳ�?*VF"X'��*<�p��ϳ�>{�09���HY�<D��f?߁���/�A��.��'��Y�sCK;����#<x���I\���?f��%a�!��τm���	�D��aGP�x����y�(D�
t�u6,�΅�����%��%~�͡��ߙ�&Sp���P�4͏��<>rI{�%�-աkj>�0�`A.�3���K��	�W��jq�I�g�l"��!�	���Mk�9��*M>�Ƙ�hm/J/�}ݎ�.o#�k�aڢ�۶�B����^>�ŬUT>1-<mAE:�ng�xϩ?�Pe�T��k�!(W�=�ryC�{�8� �)W���]{�$��� �~4�3i#��y��B���A�lC5�[�ƫЪ��Iԁk@�����$�ܿ�^�}�T���������~�eHw�FKEm ۻ,���w���#)З�*}��A)r�L�4�v�U0lWl��jvq"
^I��"��[%�;���b%���e��Џ��d|-���II�t����+
a�<^�8������g1�NI(�j&�����"�ڸ��{jƤ�������� |l���ۇWs���ȳt���"���������>����ؚ�D~�|F����=y�v챡:�e�����Z�x9g�3�{�TE�pH��z��,�瘲��I��ځ�v~jq9u�D�h�ƣʻU�s9����?�K ��u������Q������� �c�"! 6��'�sq��[��W�m� U'/��T��̮�U	@G�J6V#<�K�Ε�{�'�١��8�'i�ʎ�#G5-���ߩI n�m�p`�{	3����300�=�xl��6��ZS�QSNO�Lr���ʺ������ߗ�VI�ȭD%�;(�F��O�f��-��A���ikkq6
&c-:�(�����T`h�KP�}�����h�c˰�m� �/�D<+�8����6�
�v����JC\J��ʡ�D�1y�>U�uy���i�PI�_R�Gq�Ύ�-/�7�a���e�I����h�*XՇ����@�F�4���7d]-[�/�{`��I�Z�0�a��I.�m�-�_���j�?QZ���n˧�3�.8�B�����ݷ�����:Ca��8#�aD�Io`\�	�]��S�(o-JI�]�$g:�g4�?v�"��i@�4P��4�6���?�p���{3v�Ϥ��a�J���t�P���&`!@T�e����jcf�qV��e>@^"%�	ֽ
�FȒ��hi�*e
k;��=���� �f�x,�����T
����j�g_K>��eᝀP$bT�R�H����3��I�k��Vw�yh�t巪��2:#)�i�t�Mc�f�?L��O��G��0!F���E�Iz�3O/�N���ئ�L�����笅$cĥ��rY�8&�d���}�31vHM�Y'}��ՍI���w,cr�uo�A��/2{�zr��2�9/��l�E�GP`��||�2���g�c4����,�`��2��ff��Tը��Oz�mY�R���{���f�f�f�B�Y[R��Z��BfڋW���;�(ГgV�Wł��{R�b"�]��bl�W��ӌ&�ͭ�d��?�$�e�;Pt*�����j+g*�m�˜�Nh])��o2�|���V9��@��q�[��b<��I\(aʘbQ�l��Bhfq�V�@?�Z�U�+�9�~G�hz}	��<��-��� #�P�B�bD�ەL�N��_�'�1B,al�M�GJ@a82�����ELX���ۤ)LI/}Ƌ�S�.����IYT�䖗��4u��"%C��|�
���)�6$O0��|�N�{�̓��	zb ����c|V����a�I;�V)�법�I~ǐ>�G]�m=Ոٕ�lPe�>w�3���X2H�.p�Eф��D�ΏK�Ը�3�G�l�Z��&���`���(�����9��$7���p4pz�)v��P���'����A��2U$��d�n���k�K!r���s~�����zP���4�L�|
1*YBE �yZ���C%���z¬���<��ȶ)��z��q���-� ��j/�TA�;]�%y���H��߱�v��6N�T9�����STF�O�m�x�I�HVma�����#��]��$��1yǯ'��o#�;�H�ɵ��+ ���[�l�Ov�?Lz]��X-�\>���Af��^������o%����
����"�P�������s朏�4a�ѵ��1a<�m\���D������ISvy ɠ����RĊ<��FжD�*�F�Sf�K�aUHa(�O��܉G̑�P@���Q��87ҾPI#����#" s��tb��T�
N.�yt|g����<���5��Q�5Pₘ
"�G �e	��(�Gu%����mpJ��MIֹL�G�m�S�ù����<\��5���B�h*^�c|/���!|���|��
砑B$d��?LX�vO����y��&hF{�R�X��;Ł�F ��Đ
lX ���M߸5[���E�B���&(N�=_�K;S��d�-�r%WI�1�rIt��x���N.��8��:a�qi��qCd����8_2B��&���Ak}_|b�����=kr���Ȗ��M��K �4��y���$+��q���J���F�o�w�e�X-�0�!zu�<�ծe���_��J*�~X_�pI|%=�q�g"-{ �ЖX`¹�R\1�R7��5�0���QW�4Z�<F��a��{@	a�-͸�4�|��e-�[0�G����h��1�2��y��'\��A���_P?�`���[�7�~��5�g���2Z~��3����o[~I���	5{�!3N�����쉏mZ;�St36������&3ɢ�aM�9�Y@���,֤7����dD�a"�|��t���c��������7ʲW��Ic��SD�{�=J�Q�I	���pE*����}�bE�����:yr;��S�@a)K��W4���P��r^q� y���}(�l��'%�~������*2CK�6u�R��� s'v<��{U`A���T'���KT�I�}��
�[~�k�<d��<2}�P��+�@���J�������k�I��{=�և� �hjOY������>!._�o���?�����n=���8cRK(�؟:��s7O�N��'�ݷ�~��n�hi���M�V���0s@C���I����p,ޮ������>��̀�Ԅ�M���p�z��#��ɞK�Yrs�b�M�S7Qa�6����͖�s�Z�_�L���a�F��GP+�����y�Ԍ��@�E���6�A{Q��̇���&e�BHL��PU;��Nb�}.6��ԓ��e&R6��"D��&Wy��?�V��$��W0��h{�D�?av1"� �Ҙ`�VRWxo�\Z�m��XT5t�/�S�3v1?>�Ӗjz"@~�.Ȇ�;.��o���+�,@�eb�FQr�|݀�EmU�4|�v���N)�V��W X|��Wq��m�l� b��HP�� ���b�X�iûm(�u�]�b����|M/�_�����!�N:PJ�@z�2T���� LJ>�1	�p�#��Dx�|�R��5SYo���ڔP�)��lD�(}YYy]��Lz��u�: �a������}�L�!	��P�95݁����e�  ����6WF��u���bb�P\��a��Pq	������VB'}�sk�u�u��ؔ�6QG��I��&��x��+��L�D�5䃰��A������l�M��u?<ɝ"�jфߵQ��Ȱ�`T�X�R�)5g�-�p;|i�ҩ�$�Ր��#�|LS���@�v�h&���&M椫ETR遷+4;u�bPي6܏�(l���H�B��	��N�� ')\c�ֈ\����a"
��?�<�MI�G���{���������B���A�1A�]�M/|D���s�k��N&��G{� ��m�r�jIW��˘�'�0�/3�����2��7�����?#�%|Q~W�ϒ�5��E�J�8KgPA=!�`ZG|�1"�~a��;�І������b~�lÓ���^���he �6W��]X}�&�:����ۥw�6{������h��������~�Z��km��s��:�E��%�*�s_�\i#0	=>1c�G�"[�9�q�!yi��{����1|C����[?O�-�#"�sOU�5���'%ݙ��?bxЇ�"Y�,��=�/��% oZ�_I��#-q�JVJ{�_�Ԥ�e�2<�VJ�kw�[�	�kG��3sc�ϮX��n����{�W�@��[r��)�Ѳ$��:묎Ԝ��މr�lj�������[1k�zl<�pk�D�n�;O��mbO�Le(���G*����źґ@���,kY~��8(g�ߺ��T"�R
��l.�D�`���	4,�� ��8�S�<��ŧ�`u-G�EyH/J�kV҈o�� ��=�0#nX���u��bj��0�����1���3J�4)��?"w]�ڕ9̟��S���#���&p������KW<!G��ab^\�gz����Q(seQ�50LKI���D����U��*���zY�aX0�d~ѻk\q�Zvr�	�|GGS&�����)9��x4��4�0��o��AA0ejxj-���m��L����T��6�z8?�~~��m.�!�=X����E�a�L�=\`uN�{xk�<)�_4:~҉^+�:��y#�Φ�D$�U~SAt�_�J%� H�<-w2̶�ج��0��[��x�����}����˱��lΞ��(7��P.Vg
W]��ܽ�7��c<5vn���)j�#[��(}���&��x������Wp�������Z-q������I����p��(�|�mA��7�<�(���l��������%�����N[�Y덏�����L���ȇ9�;)Y�$Ŗ|�Z?��jh���X2��ƁfK��m��3{�oyq���e���Ru G�/�H~!7�݈��T|+�b�v��ū��WVc������6j�T��AaZ���9-?�Z��)Y8/��kJm�\a���-(��n0��;��nc���XT���Uj�80��9��L�W�"N�C�[(Fh����v�>;��Q+"��*�������j+�g�ul��f��^߶���
�_���]pM3Y�^��������ӿ`Q*MSo�D��4���y��PǬ�9�#� 	4����L�t��f.2SR]yHI�z�}�ĥmF'#0E�Νݙ5.�	��q�������_m�[�iIY���0��%ގ:}�
�Olzݮܹ��g(O�;�ʪ��:�%g�2��t&�C'���a]ӣ�'b�K�$cr���އG�S6P=GR�³��Y�C*�5������H�D�FR4j��E�l_RXH���q�A�W�<��	Y�zkL��P�B��]D���)�1 �0�?wq�pL��À*�ft8z�ӌy�_F�v0�A�,G��%��9>�>��EO�f�E�Lw�}���?i��5�/�}����Jq�Y6�A��P��g1��7��~����~9�$7��ї��ȧ���7J������}-Vi�v�����p~5c�}	��c^�� �kg7�'DA3��~�&.�н3�pY�����%��R���Sţ�InA�ޞ���h�������jÙ��������F�oI���jtJ$U�ͫ�a�A#�Nk�7���y'�YRz�x�T
���	p!g��}�m�C��g�6aَ���wR(�$f��ϟW�2;�����%n逡vJ$i�Q�k09�ʾ%��)��_�K��+4��ED��n��H*���	�X�$(���0MZln��](�N�������Ӏ\'��H[��rQ�1 G�-���$�%?r���<d�l����N�����<��;�	���f����2�CNe,f
�c!~=7��١�D��󝳌�?}��8���"w��սE CfIm��n`k��	~�h?t<�z�S�u_ �@�"F��	���
��e��ꄂ��A�vu����g��]DsV�r\��#�#��J��-�������i2��Qs�����zA����.\Py�2ӫ+H�PT9C�o�sya�XO���	֊I���V���ߩ����2	�����-�V1�'�GS�h^��Œ#0��4�^�4N�=�����K`���t���/)�&�=��ٍ��i�������қ!"��I�*
�m�����N��.B�k.�ux�ǹl����w��)LjZ�Tcy[�����q�z���1�NW!����h�����)��%��*0��CQ�����'�����@|��tJ&ҫ9�Xrڛ䗓�6��B�	s|���X9�y�b���X$u�~��s�Q|b�ɲ֕�=�pڔ�.(� ���t*?;��$�+=Ө!܏�k�+��#DUt�U���+.�NC���y�J: k;�"�.A�����=G��{}�x�HCρ���Q	qM��3]�=�{���z���y���� Ղ4x�snE/�pDVJ4a��,[90I��� �0���MhL�x5 h�(��q�>��Bb��e+�k���=���D��$��>�G#`J9��0L��`�xY>�3���SBղ>}Ѥ8���&�82���=�G�}�ꎵ��8�L]�	���ɜ�c����69�	��-ග̖+�`07���deɾ���D�1$c���+O���t9$ �g�Z��2�H!u����!W�y��*�i&O|�����D!bB�CT�E�6C�!���XC�a��HxMX��~Z6Ǖ��5��;?��;�کu��e��-� a��o�A�kV)	m'Oq�\j�e �n"��-V~"����	�y�����_z"��������!>a'�obAnr��L^�yO���l�o�G)p����Qy�b��c".��@���v}�X�M�l�
nl��P\��c�(T��Ɉg�����<:�P��w��%�ׅ3j|f�!|�L孕�
�'�R��w����߿�&��FN������DP7O�6h�A�~&0a��hU݆z���*�g�6)�I3c��H�GY�����{�HQXX����ѱۜ������꣚M{So6L68�.���T��ɅR��k���0DU^����ω�r*l�u���� �O��˩����~�ż}�\��d��:?�lu���N��-�)�I��q�SX{.6�������ގF�Uk~oŌ7�/X�i^Z�$q&hO�����)���z��9�=���U�#�x=�����K��A�-�?xA��f10�r!���)@��F_e������p��M�gr@@�.X�a3�I��úa3���dw�:o�؋�Z�30��ꮥ5w��V�,�����"�';"2�#�|�=V��%S9�!㸖��]p��'Zb�F�5t�,��a�K�c��M�S/��>ԃ@�(AjN\�����3��Q�	�A�R�rD|j)���K���.ɭ�[�!��g��\�pc�{>pݲ͏a�rk)9(�t}	�s~���*&����_�X��e'��a�s�t�~RX}���-[뷡�^���I��˝p�D�{�{z̄@��b�x��_Ҵ/��b@����> 7��C�r)ME�
��K��م8��\3҇�u
�ei��
�@w#�Hq{.��H�A�SCuj��0�(o��d�_��5;����D0�9�<..6`=Sl���F�󠽁r����򭩴��iգ��.�j�:��&Z�,Cqe�y0F�~I+4����0�8Ү��8J\�<jV�KÅV��8n���wBA�s�x@�rQ���^��ww?�!<�:]�����ǆ~�i���T�$�k�&fm��H������Cɿ�͔���G�H�{�w�c�<�T�]�[��{ǫnyzO}\N%G��*�FZ�x"̒F�b���w��.�����4�H|Xug��y����1�ظ"z�e�;���p��PQ�1����4�I,%��xa�����hR2���*|9��g�(�	A���?��5�D������K��5#��i�]�����%�L�����u�����7�=��B_T�n�Hd}EV�*��U��9'�5ץ��]�"=�M����f����)fN}��q��e�����B�̱��D�yt���5a���WTcbWqU�g�����qی X.�����[�l �Jo�wWq�-��}��x�{�+z�f�d��:���@�).d��6��o�w��JV�QP�k>��l�x� ��?I,���I�.rV=>�h�)�Ͽ�_<_ƜC"gr��r��X��ZW��۽y tP��sP�Z<H��{Q!u����"'U��ai�J��VL	���H�Q<%�E]ζ�$6oؙ�o�m<�n �l�>�v�3ʠ�˨~u���g��ѫ2�����#~���l�!� rd��ZM 0�&A�X����.�����d������@V�ڀ�����<]��'k�5n��#ͦz\`T��	N�(��4��ϯ���~B0?��n'�m�|\L6 I���MuP�bF���v-� K���63��m4��r���?󝽳D�E���ql�G1��L����w1��X)���r����Q�qG�L1���$/���������DBKEp޻�q������7��2�N�:+n�e�XhF�� E*$��j�X<t��:��Ӏ���]��vvq��I~N�USNM�E~K�NN�"J��=�@�@�T��NF,���))}/ofGof��j����4X?ˌ�:��=Os��KX}���C������;\V�)�30��n�3��:�"���Z�3��Jf�Wja���@б��.,����#Ӄ��9
�3��O���+}[�|�r�O�{�<|O�'������&����5]�m�<側Q��!����=(9H���2��H4B�
^sW\����9^�)��՜��KP~m��`�W�}���''�L��<Y�VF�V ��ٜ�o��=��s�,ڋ�t�ν�cDz��^��~��K�<��9���SgO���z13�3>��)L9�"]�\b��V A���B�Ϋ�S��D���K�w�E�y2���NF� ��?��U:����.�+p�P��a����i�C����Ɯ�T	!�|�}��|n���-n:`M`s ��-�+s�:Nr�_�����^�53�X~��. ��q���U�{�9�FA^4�ٹ�Y���}zӉC�R�L�Ċ�﫷��^o�i#�rb��@�B��aҶ7���]7�PKu���>�� ��i={w�μ]I>N�$x�>L��|�W���w�����4.G��������,���h�U£s��t���}��*��[�y�gk�N���^jd��N�ƶ�o_�7��x[$��Jmȅ^jyc}f�,o��)Q&^��х��B����0�7�R4�܈$�Ԛz'��ɢ{H��tB���6�E�L1M�焨x6X��*Du���/��&�R@�D��ڮ��aOHb�dcV�P%¥�Bm�S;�Wݵ��E��𫄋:�q$���-=T> ,�u�� X��}����m�����/���.o�?2��	�76��p�B3��ŧ<V�/�_����7.b���K?�b��#<�	�6��V��-�D���ۅ�6v�O�E?@��t;W�:k�����̠4L��<��+���7y�\V��tf�)%�́�7�Bۡ�<�d���)��?�+��|�묈7|$31�|�'ߴp�A+�����3d\FӰ�["�/{�x���q���P.֊�
�v�x.��K�F�1�X�P����hW�Ca��D/��F�|/��;�r��S�;֙w˺!�K)�k���Qӂ?�]�ϰ����FO�7c��A;B�g��@r�.��� �\5�zޔ`r��Ŕ"���bBtr��Q^�?�LE�b7��9��Qu@���T�m�=pڲ>���RG��H.8�^���1߀K#:k�K�,��W�줖�����x�$�N1ы[�N�[Ӕ?	8�iK�2Z�房$�#����E1'1�v��vq��b4+�i�+�W�c�qB%�09�_p.A�
	�����ҏ+p�� �j2}r�� �tY��G��{d�;pc"��0��<���\�x����>�)w! �^1�W��t�\�k<4�X\�&<�h'KBz?��=����C@)�����-��}�:�|�/T�o]c��'�n��
n���Ҋ����āܖ�)F��cc'�:������<��a�'�KU� "��çyv;�1ƹ`�5b�J<�gqY-P>�\�Tb�&��'�<��/	��|����|��;A���~���gLU��yc�;K2y0
��y�b�����,�W�t����2D��3�����'��%��Q<�M��,�\�P�b���㬓ʍ�6k�I�KA���l��>�F�Yf��[� �TLAl�����g��i?~���6ݫWq������	���5B��(E5�W�wj�Fz��t�sE�8��s�i{ת�V�^���j�SJQ�߷�4u�"˲�w���:s�u��# jl�	�@�8ylbǛ��D��!��il�"��iȧ�c�1���O�i�/L��㓚'��e�s0t�,���!U���N潽V����{��yy�
�y_JDu�M�w۪���7�{��푮/��uuQu_���)��|�\SMf X���nO�8�֌6�e��/��x�|�������i(�J;z)��	�����t&�<+8u��0�y K?�ն�ta.6EM+p`�Y�E����lp�$o������S8��Pp�h�������[~��e���iA>?��2����BT�t�8��(z-	�+�ʲ� ׺��X[��z�z��챽|�J��7�FV!�w��t
�wV8�9�(#�k��AS"�]�d��n�����|�l
w<c�՘!�Uzm��^ͷ�!�J)OI(�ޢ6����:Q�w��b�I;+&�H$�������Q����D����o����x0D�}�bd�Ą��Z0��=l���y��R���U�פI�:���I�ww����O�'�X˷�v�WN+����=+��[�Y1���;X�ѽ2C]�w��6d��I(� ܈�D,:Zw��b}x�"3�8��}��/�A��!ƝDMl�]�0��s�+R�[y�XN2��9�.�˗�5.hZ����g��j��V@t�Y�{6�����YA��b6�Ґ	�6����&�<���B����}�2�V��c��������#�m�."���7c�vOt)�@ �7,�]�q��N�Ǐ-��޹ʇs8x����*yt]�b��M�C+��x��k��J�6Z86x���*0YC�s��VJEe��LKfn��ϥw>=�}N������]�m>w�j�<Y��׶٪��,��F8��V n���:���F��>s$��t�x|UG�y�x��(-����.�6���#.����}gg�iGr�]G��F; �y
�-����kއ�ď��O��i�^�sf�.��͐ޠ�W��Wo�Xn��}�.�j^�����&��ͫ�j&^r�s��dFi�5H��C5A��^�GO���/��wmT���(��H�7������3R�Օ��Ŵ��*�~vv>�q���J'�f�"�.�Y'�fǱ�ax"h�G�Ax��*���.s Q�Zα���Dq�(��7r��;H��'O!�_��$�K��+F�Qn�l+Vv{�[���F�o��JQiq�{I+�6�]$�B�yS�Mq�kzv���;�t@�u<��0	�o��B1z����U5_"�ʰZU�
4\��Vܜ{5hd{�`76�	���4qץ��x�=+c�}NN�V��'�_�H�:�abAKj�!����wK��R���|Ba�X��C]S�"Z���
5�`�e�L7`9m�]kظ[�p)%z`�4�	hXL�M�_�
Y���VSs@��>@xR4�-*���������6>�f@s|��.����H���Q�OrϿ����@��`/��	}e \��)Y>�$��V����y!N���v��I�a�h��'7�����g����ZxI���p�P�e��J�G��j�ڽg���~ iDԎ)�/4=44�ߎn�B��'wl�`/�D�R��X��~���=�15�⟶dmj���`�T��y�Z/�>�=�စ�j�>q^&I�
Q���\h�S�R�qH��LCz�45%�����rC<2�`۵{U5Ћ��������J�/������Y �%��2��8��?i�B������Ϊ�h�K�L:[��)
��I����a�ظ�Y(�ޟF0)�<��!�$!�>ꉡw�V�g�wE���F
; MY�e�=>���KD�M�\*���'i�����A�����\OaQ�j�i�CP��c^-��i��D� �D���L�w6�jo����j�����^-��Y�@��{*�(�*���p��n��F<�:= {�9��t5Qv�=m�V��U���:�̣�|�o�ʃ+[]N� �q]]��ݸ-Y�L
F1N	�i�И�[�jL�y�a�1鋽o<��k#�UA+/��8���;GF�r'����r��3�pQ�/J����;,X'��?�يjX3TTm�5�j�#ĶVL��Zo� �sk鰑���/%R������5�/�|����qC?(�?�,�{����TC�\��=_�Pd��Gp��T���ܑ���}���!K��+��$�,-/%r�S���
�A����B|�k)7�����棇`��Q���%�u�Dl1�q}�4t�{{_��F;��-(���$-�pW`���6�~�8,��@�b]�"�L�4��3��C�'#wJ�7�N�q������V��w�gI�ه��Hy#�J?K�鄁���U���jH,�L��|�QBK�BTn�^B�*�||���UA���Q�rwn�@&?x3,�nl�|�	�XDZ�A��W~o���?����E0P�ɖ��Hyv�Q0�����ݾ�����j�ĥB�GU��&���[�!��k������3�a��nu6�&/`'�1��N�|W�emP��J�L��:h{¥����M}���/W�bD�h(ˮ�>���5�Ps�b�����6�cȥ�l��YD�	���G`p!��b:��@�H���������X5YCd��&���w�љNi�����p��)ؤ��i=���:pM ���sD�mng^;VB0��)��&�T��Mi�Rkk�i�x�+ë��N�O
����R�',�->�;�Y�HaO�Bn�r,�F�H�����'��N������q,�>�����@��lX	�o�,u��9�:��
�K�_�����A*m: ���d�{�mo��湢����=߳����tJ���RHrf �͏p3�r3��&Ǔnm��%n��:O�U�7�t�#��g� M�L�Ĕ�X��	�ژ����(u����fb3-�N���gyIdsn�q͍�.:���=&�#q����t7uΕT(QL�P\�
g���%7�|Y�����&'Q�N}��-�6K���(X���!_��}y؅-�vqoi�*��0��=`G���>'��	��0��+��<]p��W��o��Mj���D>�=�U."�ko.����y}�y�y8����~*���w�|)�\F����u��yA���Ջ�E��a)���uBQ&����W�����&-��qF��m�Itm�F����p��Ew!�{V�/2�W�"��dK�ª��{ݎmh��(�:ڳ�J)���O�F��W)�x�x|�0�/���ٙ�s��ȱ��S��0��
�Mfb6�f�&0Cv�"�𤈴�Ԓಎg9o�ɝ2{*��L�ѳ�Ci�!4�����}w�������]t**��]��c��5~h��D�Tƣ���Ah���2��s+�`�1I�/i���@
��ߵ��03N��+�jrKAX�ڭZ�w�SX���B����j|�s��q͐'�>2��xM�R��_�G���6Wǃ�.6�Ƴ�L�`B:�k�K�F�E�3��18��?����;�C��úIX�8*G��i��H�d��c��B�~L��"�4�������De�[�K2'��)���>+ ���|a���>�-~9�y�0%����}G��݂z����	Ho�O�ҥ�?n�E�A\��{H�<aC��W��3\?�!�eҲ"�ꟶ�1��Y��Bs��	�!Nvu����� b'��V�H��ql�!���7>Ati]�ub*Z�/���p��Ÿ`꒍Aa�ɤ�\^Л_V�g\ݎ9������Lq�h���1<'�CD�\YOK���Z�' A�[� ���㉷풬��b�=�4G��Y��z@�^�0MC�k�^ayvs�+N��ì9�ʹ�7�pdo��^X��V�<r��Ž�t#�J5)�Q�w��o�7/�;���1N����f.�e�r:��`NŮ�k����=�;�D Ht2�y օ���2&��&Hc̎i��l��W�d�_}9�b�蔇���J�R����XB(��KVa��|bAݲ����[��co;�j|6�&K�g㤤�#o���m���\>�WzLp�^
�v�S��i�J��'��K��/�"��0G�:�2�Ȃı��`��a��2��5Q�)�pl=����Y�@k�j����8��Ӄ%��^��>q�)������v�T+�G��5��S�i��\�1q���M���"�-�x"<��� �~jeP)���_l�%%������62�~ۥ8|���c�vI�@�i�IT�C!�ժH5.��cV�� ��H��<j�i4���*��,x�|���2yo*����:��m�:$�=�~�5���I���7l	3�<�0RK����s���p���x�~112��U���*;���߭��� >X8sR�����^$����x�H�2q��������y�6F>���������ō?K��A���c`��3��w�M���Y�n6�_��դQ���<�syZ��W/�xr���g{Z_gΩ���i
��f�$	f��q�_�z��M7�����6%Țy.��@�7����O�e"Ӡ~��x���5�|���O�G���"?Y�p��U��,L%��2z80I/uQ�������onIvb��gu��%c�*�Z!��+C����i�3�zE����)�����Ab��$�z T�=���U�(�<���s*�a����6-�*g|��y����d�X�f_�����U�O�� , t�SF#���?�����������;#��H<KQx8��V�]r@�uN� P8� =|�ڽ�!�n�0�;(��G���q"i �JK?IU��
+�ݯ�\¸���p�j�;��oؔ�M���d�H�7_y�:����E����	kCq��|t��_�j��=^�=>�d	�Oj�C/4�p��ԋ
 $k��������Ɓ.0BNd֌�v�S��݂C�/�xc���h���{�Y�!�4:�`m�óe;@�l0cpj�,a��R�Q6���ܶ� ��!�9O�� ��oo�A*h
�����9E�u�H��B˂5pL�B�X�YJYL� ��Uj�*1�@�c����Z���\uI���yo!c���G)�?��W{��N��:�M�1��g6�§�ᴑ32�K0��,��3��V7��7-��vƴg_w�����G_��ت�j��	՜���i��%d����K����:-A2j��x���@I�N�0L�5�5������u[�J�Uɭ�J����Wk)~�25�x�B�i6�y�9-�#���\�Z�ǿ��7it�s�a#4v�"[��ئ<cӌ� ���@�H��82o��"x)ZC�?���\����.,j�B��֙J�[`������6��舓i4w�:�"�%��X�:*�a��ޑm�v-K�-mEQ�Q�h�J�A��s�{ο¿9��Hȴ�
�U�g���=��)C��w������S����U�{3�"	��]?�J�u�>�
��>���@3�	�_�;���n�.��?=݂ҏ���4"TB�6
���K��3�a� w�g��ڭB87�� x���9��#���SA(��l���0�o1{��,�\��O�i*�z�� ��TԘLp����5]��$.*H��&|ک#B)R�h�.�&U�A�Z�@؉e��Q��;��/��X�>�8���>6t��Xl�Vb�I��'��م<������ !7��L�"��a�(8���
v9Ј�L��M�-��+�6���.��
!Fa���4\�h���Y��H>�*ׅ�6�b�|ܢ;v� �x�ؙ��$��)|�5���ÑNԒ&!��}ǆӁ��tg�Շ�s�l�>�h�`J���K}
U�8��&�z<�,꾦���R}�i���_�Z������[���8�J��u\R�xT�?�F����X��pxqڇ�qU�?,��Z���f��f0�<7͌ŷ�Bh��뻕�<GU�2	�i���$����ِ <z aԆR��S������w��T$�bc�"�x��c4aM.vZ���/hr�����͹(n+�|���i���#�W|���J��P~��)C��w�\��lv��GD/�4����㑆نH���A>HiU�~Nd�nk�\L���g�Faf04p�h%�� �f�D�$��y�:M�
�+�����a5�pGO=r���s���a2��T��8��܈�I�r�&����	\�D�ĂK��v7��r�㑊�k�&=O0�l{B���1��)etKTU�,j����q1�Y�
�h��d�1�	d�j"󅋗�h/yp�/2�r�ON�/�9?�u^>I���o�#x$�l�7�����]�&C.�wY���i����}Sz���b���m�<�4�6Ud�f��=�}��8PU�P|��!Uc��"������L�be��k�g�	�������/S0|t�Rڏ5���n��F&0�	b�Qؔ�]����C-,A/��5��&�������:#Kx�/�ݚʽC�#�iV��ld�P^����m�Rj\w!��To.�h�<�F ܭ�6.:W>vG>0R�D���̓Im�>��;w �c�5$%�6av�ёNZ����k�Nc�9J?m"��#
 ����u��O�^�ݛ�����%������@�n<|�b�2`,�N�t5!H���1�&1�(q�������L�Sγ:%��R�%5���z��`,��^hjM�@Q&9�ruf�)��X����W��<���Ӗ��w2^,i���!�����ݻm���;r�i23yg�$��\�Yy5�Z����ɥ����m�4�OcMI/)�[�j�؁����M�V7��e�J<��ZOmE26u�6y�J�o�,�d�fK{�ǀ�&F�y��-���I���X����{�sI%�з�(<b*��-���Mu�x���02�͝_��9O�y&�2bg�����t��V�ˆB�A$"�T��}S�28{\�5�4�r�֮L_��i�-�?P�E@�,��cFN�Umu�8����	�ȒJ�u��b_}�o�q��ݜ�5,ue�[��Z[v�k�, 7�Y �i@쮔  ��`�?�B��݉���	��)�mĿO���P���c��[;�DA��{�qG�W�Ɵ�@��~�O�s�6o�a��gq۪O@�Z��>&iQR���+`N��$;F�O�d,����ԋ�8¬;ip����S���!���r��+�"l����$ ��&+ooC�\�2��0S�	we74b�E�U�h�Ul@�egΎ&h=<,���ϣ׺U.���o��{:\j��}[�Q�t6����IlS:�JI[)����l����C�Y�����y=���W����P�ȍJB�Ϣ��aA	�zUe-/��ξN �:C����g����~�6Ux����ӯW�w������B�*��L_�D���<�e�D�����l���8��Y�U�܄�}ͦs���5ad��)��3�z�mT�9�c�5~ᒹBYQ�[��{ 5M����Xj������h�5[m�o�#<�L��Q��f��A2f�@c~�v��vY"�|��y��.�Ⱥ�s�3eX��f��*���}�V>eV�4L�H[:�UX��_�ϺM���+�}z�����ān�?'���Pc�vݹ�����/�i1X��5N�rS�S�\����PPm�ѵ��,+�oS�)[�M]Ī�w���~ �u�a�w �*�O?>q)lz&�����(�r�@A�WJ�X��?�)r��%������B�+k��]?����S&�/��1���]u�@`��ӽD��`ΐ��'(5�6�����5v��ՙ��<[�>@G��j�#%�t�ʺ�H���&����Ir]��Ԍ�鸮�Ĺ�6�C�v�Z�F�TM��������uю]������oԾ ��@Q�q�"�#s�����+�0�j9���Sk����o=yS<&��|*�6�Y�<:qu:F(B�W
w���S&��t�Bl�@�$��=cu��$1��L1&�B�'�`](\$��)� �r(Qe���4�
� ��З\Ck F�h��9�f!F��r@D��Y�8�l�^y���0����L���j��qǣ�w�O
�on�Cb�#��F,1�0`�a�%jӀ[��9�X9���>�7O��H`~�7
b�\Z2���#R*�P�3*���rI[|��
G��K`}�<�htR� �Q�9��9R�J]�Hx�#ގ�$Cn�C"Ĝ��|N�mO��mԔ�Dn���@k�H!�
L�i�tґ�y���R����	�C$L�hKJC~�-�--�|�������>��8�oy��'V�����y亡�l�1Y���P:m��d�	��|	��8<���$��W$;0O�uG�D���+����� A5���G���TA	��^N�O���k�L��#A�
�ᝯ��}$�����nQ�Kj��#���D�P�;����q\���kZ3����D����Y��#I��P	I>�Xx����%`�	���a�h�Ɛg�V4��l����.��j׹��N�z&����N�넊_z���kw��$#�����ݻ�4riD�8�� �F&����=����@5����X@:�,#��E��?,V��k��������6�N�=հø�K�쑜o3�]�D F�U�C��)�ޡ��2� �ma4%�;��@,r4�B�b�����bP�THl��PG�!v�d?y�h�&��ۦ�����v.QXR���:���Eķ�Dsy�|,l@IЪ�CmE�:ժMϠ�<��)u.1{LQ����ۙ�YbhҫL��t��1��u�\1�GPO'8gn���'
#�7�����+$n�w���}�Ǵ_2�+h�%��F��&�{�!�� ��Fh���_��"yY��[Sژ.xHew��{�8<�e:>W��񽔍�x��G���]������Q�y���HY�9��0] ��زi.X!�\3�c��N0����[(i!���y����.�BФ�쉖�oZp��׻~WE�.6]���:�J1�"w�k.������4�(s��#��8+����}R���KR�/��bS_��(n3#=���c!��A�Ro�lVr�yR���]br|�3w�@��M�c�cKB��=��j��"�(��,�x��*麒8~v�=���H�G���[-��!(�j�`�`YolF7k!�`	�P��xq��X��3�f
;���8�7�����Sn'u��Vy|���J&6��
A��������֍�çv�]��F�����Dt>w�@���]�Sg��D��}O�~`���{{� 2si�ƪ���=>��C��`<����w�8iTD#��2�#b%�$>9uf��d��������@�-�HM"���]9��L�W,a��HQk�x:;n�c?�<��-�T�)Z���;�\�5��$]*�����/Y�i{����-��ݪJ�Ĉ�pU����p�58y�`���^Y���O
�6�>/��l�'r���]�
eP@��݀�o�"+����.t�ґ.f�֡�~"��3�n� 摜�#��P��f�aʱ�.^�D�eUb�� ���1���1R(q	��3��/eP^T+�:�>LwC6<74�)����F�㝩,.�?������=�Y�1��U�)�Z.��G��ձU�xo2�����k�"�O�,=KwH���,��Q�F�z.=�b;,rr�}'9�+��D�kM�VKz\�1���R1��Buq�إ9�	βw�lR��R����(�e8)�Z����K��`d���+\���d1��xpZ0��SH��KޙUT��u���(Y�Kd�>B�e���;�f���<d���:b7�e��ݠ����ǣ�J����_G��U��Z>��`|:.����k�Լ��zFVIT��넴8f<78o*��3Dʁ����2�~��%����J�<������������QtϹ�?fݧA�����	 &�A�t4��5����"��+Lo��s2��w�S�l�x=j�%��P��Gۏ)�g�8&�V�� &Y����*H�ޫ� ?�0�OǸ�,q�rS�A8�w|R�qN���A���g���=��,Z�J�L&|Y/��F���O�~:l�犇BQ�����\�}<���������on`�/[J;�Ouhq�'��ؔ���d�h��?�Qf?'�Q�L�~]|�L�e�ϼO�����ޝ��&�o���â��0,
� �W�wk�2�E��V���U�Ѷ.a��K�f1LS��{EPy�5�+m,�"������m-_*�Z��΍Cپ�W�۾���	ؾ�`z$��l ������K.�9�~�"-z��r�&nfxڻ��ʌ ��¢K�KuM�j��75*ak��`4�W�쏸�f��R�&B[J�˕5�۸�a/�f�/8�Gb%--^�w�����d�9c|/KQ�C���`�(�������[ZCEʦG �Z���!F]�.T�X���5�s׀���=���i�.(V�('2�lS�Uh�@�}��D�#�s9k�j���XI<��D�؞��{�t��<�S��ZȉQm��)��Y5G��)*I��Q��qZ4��xy��m�q@���W�ū:T����褽v�=(�ul�A�er��al�5��Ϲ���O3�zT�����M���D
�)X+!i��1_#�Kqr��洇:F���ղ��f˾�k��PMb;���~�L�M�.j�xz�vH����bY�������Ͷ��5��t�ވ���7��(�fǤ?�����%�A����3�JlF� �A���Ḱ�M���F<s�g
��J@�%��m� ��u8�=�F=.Y�f�\LV�y��R(S�h�6أ�c�^�sɹLzςT��a�C��C_l�ՙ+���*�����+����U�����Q�����G��ػ͒�ԝ�����.�~.������bSJ�b��X����.�T��9�5��";�>�*�ֵ��U�����%jÇ�G�rt��j��V�Pz�����E�:�3�as�����e�N�?��z:��.��������JP����+e�h���Q
oԌGoB���E����{�R�²�-8��&(�ZB���9���/f(��F:�@熚��͹�.oa��bc��+r5g��O�ԩ75	�Ԋ� 送����ܓ3�/|ޫ��6����%<��ޟ�K��L�p_!�dq����A�����#�L���[�'�[C*���$���}1o�j��Ͳ|�������w%ҫ^#�۪[�}�9�4]G��Z�/^��n�d����~�恿H�l&����r���\Š��QI�ā�pp���<�Rs��`H��|�
?�C��|m`�����D�W��=TZD��ׄC�p�����/������"��M����0�h'�G��V%��S$��}�t�2�0������m����L��hMU4uTI�<ռFP�|�K��5Zt�����X����v�8"���/#3)y\ȿ������K	�u��~L�2�� ��,.�
/�i�d�*�(~--�&k�\m+ho��-�s�q�yz���[!���-V��4�+�Wl�v�k������t��p�5�7JV6���r�x	ݽb	��x�[��WR���F����&�U�b�D ,'��l��CCF��z3m��5���{��2E,A�O^�G;�Py_�rg��
4�Id�IN�Jr����`=5�L�}7	�����G��9���~�u9��">�cJ�J���y��[u����=sM�H͝uX���7������Xh��'��Ӽ�Gdq9�M�t��j
�O�Xo���R%6��5�\G���#@[��M���w9i.��  F}�C~��� P=dm��pa1�.���i�=��W�Ɍ����Fi���G�H�l�7h���)��_�$��j|���'fM��#4w`�!��׽P5�����׋q���D������|G6�u%K,��00�yA����&uB�k=��%w�:1=�������Ow��0�����9P����Zk�b~��6�h}��^�-Pq�ѷ2���	�59i]��P?���oIV��s:Pa���hV�#q��/jI.�#��r�{��{�/��R�B�@Ι�KLo�nB��O�Nd%�k�g�ނ�,Y��j�i)X]i~�0vAO���<���9h+?C�d��0�>k�m�h�wTy��B{���"*�_8�����8wƻx���愷ϮB��A�~�!���v۠��P��6#,���e��D@�U���\�]9��>���O3Bv�wo:B]�@4��t*�i�(5�O/��d႞m�v,���,}��1��F���[B���[g�kZq������E�U��Ç��=�r	�=�����H%��w��Ҟ�i�0�xL������#?���+�͚+R\J�\:#��Z5�"�;]R�Q-,��88��f�ODX�w�V�ҡbb�_�U����ڒ29ֳ5O�T
W�S�*51��#i�5p���ˠ+��Xp�� :���@ ��A�&S@m#2-C-�%�˒��?��! aA ��F9�@"��ow����8�1��Fx�	{H5�4nT��7�&ju;tV�ש�~Iҕ��#c�.��� �h}Q�@S���^�AI�]��THL�	��hB2���h�:M2��$D�0:Y���ȏ�/pଢ଼���۾)$�t��m���w��S�I��R� ��=Пn<�M����e(�R�ܠ���}?����5�8����9����1��0Hv�&���p���(�`��b>�|H��	�kw$���b�`�B�$�x�#=�O.��/���#J����⧤���{OY�q/g����b�]w�T���T.��w{���aΪ�ِ�����F�~P`8Xk���ڊ^V���7u0��R���Nu-�,�}=��*q�� N����!�c:�/FᵬD)�mZ�k]�j�l
�+��渮5��V��d�F��H%�n��|ưh4/���A���/L������֤.�ER��BG?YOt����ҋ�2L@���H��o��b����3��}�?~����	��b�X��C���A�1���p�j�u+PΎ��k�����ǿFm(D�$�ҹ� c�M�&߬�h9��jup�/�6�C��à��M�p��?£"�[���p�@��%�o/��%t�/����væ��E4����.��L})�P�H��h�-%�p�o��[@I�^r��.Zc-@�ٶYwf���98z��x@�T��8��[��-C�� ��E��6������up
 m�������1E5�]We6��x�{5T��3ew.Ԩ�zjR
���wP!Yu7ȕښ�Tw�.`���v^е�{-���H}$�����|s�p��D`��@���0�����^n1�}�B�N�3��`b>�����u�N%�V,SU����p�����
��ЙZ��E�"��?�lx$����fBÉX�VP���F=])`!����/1��z�N���Zv]b|m�h,�Py
%p����Dw���Q6��4���W���C����~Xi]$p��o[d���v�t�B�]�2�ٖ���ܛ���5]^`�σEW���;f���b��p@{�oKaGr$�R�*�7Wl��4��j�5N�t�Q�-a�5цr�'�D�T\�/:cg���X��Va��5s1����� �Hv\<]R��޶_B���ĤN6z՚ځ����F#�q/ި����;��ނ�K�\@$8�^'
*�+��s����=�Uԥ�#A�8S=K�6�v�{Y��Qݓ��	����@\��I����:˾ܻ4�PK�c���	C�L.^?c�ʾh��W����Y�Wnp��8Sa۬=º������ni�*�#qx-׾��r->�]�}����~��9ƪq�[�3~�X������.�^~�]�[�: 1y��bP)&}w[~�1�b�%|��V��fC�RAjYᝩ,�:�~D%k�V�	NV�B�(1"������=���!��$q����G��ߪ�w|�h�p_��yN	���1�+�:��Z�cDK�X��ap���T)���"���<`�#�N�]��D���5V#�mhQ٣M^�V}�љ�j��Q'2�'I��J�N���g���*@Md�4"Qm�|�:����� yM)��I�@hs׵�i<��{C)7��9p>�3�D�l'o���j�C��;�P����!���&�)�d)'����0�bMK�k��Y0�����$�gBg�]������ڜ7͓(�,���/����1/���7@�:��z�ㆷ=���E���;���N�sR?�T|Ѣ���� ����nA%�u5�iΪΗ3'��(}w��đ���ha���G%�ȡ:�dۼo	\Q��	N�`dO������ɂ|�*>!	
v8#�6 Xn�!E�=BA7��>�^�$̄���u�0��I�~�HY7�Q�\*���q#����;���c�QA��!���抂��n���h3�˵��͗!Ce[!S�1B~��F��Oۄ	$�ʿ��Z�O��}�|�GnO�r�
�vL�Ծy���������; ��& � B'���4JH����ti��Ӝ��(�b�ք ١����^�p[n��v�ϭ���8cAy����k���&?80�Ʉ�<5�Jp��t�_Eқ~ �r�i�����V�e���J:��|FI��6x�:E� �
x7�5�))h�0���̈́y:[��LzyW�~��i�)����_yt����3��;�?�a斺�$��e�`���������_x?{#T�
�w+I���r�˙�iG���mGCo�:�i���(��A����.�v֗�6�h�'G�;�א��\��_��z�ڬn )�CΉ�}��LQ0���z.:ߥo��w��.!QԏX������
�ś��g�0�ꊺ=H3$).��#Ak����
So��˿e�a����iOҺ�+��)���!�u��"���7�g~|�hj�':V��ܙ�/���-���m	.�{�N�p�£NkT�\[T=�?�5X(J�;���cԡeO�����3hux��� /]�{��30s̪�8�V��
���P�m�>��`��k�[^����c�[}�m��#D�*��>�U.2L0|�5����� ��ɦ��\
=��1ew��]���u�mD9d�v��g#W��or�#�^Nt�����3b�=%��U��f�(MU�y��E\�䀷��oyD5NQ2�A��f��9�%��r��+�s�bv��B�ߡ���EN�d��q��F�,��^O�� ���(������{%:,q�mmcb���q�V�-_�!+#�d#����9�q�@b#�a�%)G
%
GG�^{t���;E�Xb2��a����`�Q0�����A���l��:cWo�W��Q�a6����ёڌam��4�ч ��'ͮ�ߔ��=��Jd�Y<ō��M7�;���~Q4|���\����j�2�w�]IBQ�ZI �b������Е�3�����W�\z�Z�5�o���҆;Lh��"T5b���4�62߿vJ�����K�0�z"�3���m�9FJ�&��S�y )-�ׅd���~�K�.�L�ou)����4���GDE�)Z�"M�8 B;j1%�o��B�m��{	���j�7��[��UgY���=�r쥻�}�9�,�3����v���5��Y�������L�\���먪ll���7qj�մ��:�HD��)��{��Zď�"�\Nq$�H>R'@�A�P_#ذɰ��|��]�Q������]$EG�
Tݩ[ه�D�r��
��ؒr�E�-f�p)�\Q(���	c�v��1�B-4`���E�TY�>��%K���;{���Nˈ(�h���T.�F����Z3Qlx��:�����K�������Cꈬ�0kf����1��c��t���%�G��_�S�L+��)t��˰kX�b+V>˧xի��  t^=�ޝ�lv�|�֓GaK=�� ���l����]��z�E�`���Y,ԵiNG�!8`��׬H�ʢ����0wB���-"�ý7�NE(�~�~'�	L���_�(���|����Y���a��Z�X����8�I��6e���h �M�'<�~��	�묄'#���]Xi�P�yY��qs�X��<���5�-\��n3���ڲ9Fm�h=��q��+'ƻ���n�~�"I�924�hk>v����/�In�&�#�F�u�"�i5ē��>���A"@-?Ph�� 9<W?
)�}a郚�%!/�YwX��3x����%����V�0z#a��+��8�c^� ��9d�Ǝ.!��� nGP��zp"���T=+bc��"c-�R�A"�7�kP��*��-Xd34r���Q�{�E򥩜-�&����P'��<'���?lw�k�'L�zj|��n���Vm��.��? 1s��wC#Z�P�N��@h���0�����e�0� ��k�rX@���#����"�9e�
�;wgm�}��,�
E��ot/�6I��� ��A���Z��>9z����qׄ5ӥĲ\����U�<W�Y��ށ���n7�Q��j7!|��d���p��!��'2�^��B�J,����~>�"��}'+o�㗁��!�bb*��9�dg���`M$�����2�d�F�1��L�&�	�w訸`��g->�V	���]P����D�����0v�>�,@��H�*YN�m���䐆��`����Sp�ڎ�1ŚArh�׉@�+�p�;b��,!�K�ϱY�{�ݶ���?���!:vKIf�&x���9�8rSc��H��xZ[E���x�H2�;���x�Զ�Q/F��E�Y���_3^�`��Z:�(	=�Dיd��#�L��¶=z�!#;���.$��JR`��SB����Aה\�ڽ�p��5�$cv�퓏��ۤ��/"�$'�?pq��:y�<Ƚ�AnN�����<F�a���hϨ��Ǔ?\8D��F�܋����I�ק�Jp܍����u�:�6�m��ķ��E�������,���B���C�TI�����n��ߝ>N(>VY0�j���Ė�1Ij� k�DCc�N�`�����O��{�|}��
K���=�gZM��2�N�����;�{rOv�ɠ��)��.bQA7�I=P[�-���b,T�Ńx�RP������B~^��Ѧ�נ<E���sY�/�+f+C"i�ĭ�y�E�c��2��lT�f���"����Q]0���'G��3X�}rt�UV@pLи�](k�T�#��}q�&�ӆ��r{�ڻ\����1�XݛC�/9T	?�,
=A��4�K�G�L(BX�P���I�4/����&��!�|���E��b�U7<��6����C��įq\r���(������K���絰̰�9�n�vw`�Qs���WR�F���� �%�Y��o���xX�W�9�7��7,bZ����״7~p.+f�I�������@��R:sW�M�����(��Dء����
������=�����3[���[Y�c��!fN�7�o�T|�Ї➮J�u��G���Q��T�>�E�o��x\ԕQ�}J��~���?7B-�)%�z��9��C�:c�7d�� ��� z�2�A\�It��w�����9��N8+���9�Ҷ/N�h��-K�k_7�4S�ԡ ����C�=�����5\��6��鼙�hh=4}�^+������t�[�CY���4~������,��Dr������`Y/$;�|R���X�k�<�43r�%��}.8�J���j<���5�4��jbEѷld�0m�pC�x(�U9 ����� ~��`������Fm|@�4��|���&�2]HFK����]/^y�O��0D��N�]�Q�l Z�?%��P�5�ꗖ�z���A���w�?����jᚊ��Q~�o�Yټ�A��_'2�O��B`����S���N��]YKF������ Obq��q�@��
	MZ�3��p��ն�W����X���1�/�\rؗ-V�Y����/�82|�1��bF6̿����c�I�MF��2���vBڝ�J��*��S8� \����FCě���#f���%���	�MCi�G��ķy�$0[���5��R�>:� BdT�S��,o;ӆ��v�\���B�CFMO�*��U�<\\0����h>w�ć�GU��� bѢ;�K�.�[sh�� ;ؕ6�#�(�rf,�l�_B��C'h��K��F���k+{ʦ�經�l��jA�lR>���b�D�w���=R���؃�d�� ��t͍��?pZ�T� ��>Զ��}�p�j@S�*g
/G��m�4��1	ğ��E��<mߺ6�^t2�|�>�E�!��t�w�)D�a�#ӡc��<�������,�H�*���[,�]�Rf�xfQ�zǮ#��]*q+�K{~�r�B��6��	�Nޕ�mo��hx̹����|L��OW�)���k�)/d*�_b�s៮S m��9��{�H�5e{r�_�8$�����n�~�أ�����R�/l�1�ы�hoGAC���4�T�:���\�YN�A�*NO���O^�>ڝ��~��~pJ��)<y=
Ed=�����ki~��<� ؂��X��#P�U�}�q4��5n�cI!�G��`�?����UFq�D^�v�6eW�7�9�A��R;v�����b6U˦..c:�-j윊~���Ո����Y�LW�R�;z8�����ߴߢ7Q`'{�}u�9��֎��8��N�[�F�H��tF@	��#�ֲ#���ܑCN������i�h�"����+����*�4f�ʳj�5�p�zp����CdQ�X��(?��v�2i���"�_�2��/k:掋eb�Y�3[[�����T͂�G\/$�:�rQm?��R�b�욨�v���r@�� ������Eʅ�Y��D��R�)BM�����n�/ڇT�k�A�{�W˂~�w%��dH?RH֖Ƚ��ޑox�����*�~p.�Y.���U�PvE1EM	�*d r�9"�u�]4��n�oYq��r�H3yuU+?z��N�ۢ���$��C˓����!�=��>DL%�$���e�Q�yj	�I�˾�\O��wmg�1j�	�GL���n���J\��w?\7�!+mg��C��UǋL#��S��HY׏1����*����d}�-�<�C�M��V[qp]����5�dܞ��� �?�X�woz�q�	i��?��m=L�S����H��t�k�+�*�û^s��<�q�L
�[^CA���a$;~�$��5�R@'(޻��[�cxIHX���.ab��3�"�ک������Y���˞������+����d�ǘ�|��f))�B� ǵ�& �aK�	��E��TȐ�?1�te�� �LY�+A�2�P��i�P�R����s�rz�����v`2�O�H��wv5N#d~�	��<�.��U�(Wv�D���Q�U���ޗٟ��	��B����
��J|YR~�WO���|{�(�Kfk��X�����z��#8�2Ap�iAX�P�a��G�����ϫ3�R����i3��[m x�l�@�5چ����Ƣ)�{���d$����Py�O�ak%$������G}�X�6?��I���7��_�p�)wd��%L�� W+�_�8��#n�j�������<;ɪT Y�)?�f$3E[�+��\4�	��ۂh��������-�U&_ֳ�F��#>�Σ�F�vw�G�^HD���b�q����k��5x����f��RQ��+�g��1����-n��r�Lω~�2wL#�=b]Ǣ�B���a#bvc���]7�zt��Ƶ_��;\OPX�Ã%{ָ��,q�_"������+1%�~����*Ea��[�\ˇW�|d�������<��ֶbV���u8�B���ŀ3�� �p�/q47Z,(�o'����~�}�9[!Io�m.o��#t�C�ou�Z:��hm���GS�%������B7^�OV��@����wb�t�C�bCU�u�7̻�����ֹ_����WTsJS�x	(��ѐ)�-v�x�~�ۘ8����Z�n���+I�����<'���]�f[��@���%�n��Јr\|�Z���$L�n���W�L�?Q�gZo_�BZU�}���ׁ����ʪ���2����~]���M:������h�U!F|T��dɆfZ��e��bq�XB0��2$�z�K�4�����z0X�n(��Z��A݉l��=��o���xy��r^߉4�!���qL(�X�������.u�$w�]��g{B�g�= B��LR˾0�o �������1��o�z�BЯͬʘ���l+����b���l�F�|��L�4�`��h�����F�Fk��������΂�����t�B4\SA��+D��o�r��]�e���C��Z�s���I�F�u����?� j�9�o������+ձkg�2�`��$1��`>	�(��%����5�@GM �mlpK�g2�#\�Z�A.@p(s'���K���r=�C�=���6��p��
�pi��1E?�ZK>+Wj$��!56����$�5�
����̐)c4�ˆ9�9�]��Pvv�P�t>]���4f-'�w��$��F�J����R��Tr(�0�����MU~=�>}��Ճ�ȱ
h_+�<� sP� �� ��P6��U�	[Kh��
��4t�Pb�Ǟ �4����mT�b�����^v��Y�
���=�0�#�i|-yn\�5����k�eНzJ�����{��̾V}Esc���E�8�1���L��K��!�-o�1Δ;Q�SF���~>��q/���-�K����;.93wT'Y�YCɯ�0J�H�`�zUB�[�qV6 -e���C�$����Q��/KYl>�sh�e�4:yH���U>����q�܆��g��ޝ�l	j9F~��V �#Pq��g���l\���(��bIme6�i�P�Dt��	����r��zy%䀼�k�sT�\CFi�ә�=֕�i�B�Vf��5J�/�H���~O������)�C�i*n�"�l�L��BLt���ޙr�U2�v���Ql�WFɯQT�,U�nj��9����̙RF ����䳒���z_:��k	�ʍd��X�ld6
f%�as�_��:��ի�L3���hcp ;.������}Uw�g*R);����	�Y]�^�<`����n�Nb5����Vl���i!�_�C��~���[����R/0zq���b꣢����E�_��؂�m�7�i�H�)#9#�V1B�{v3r	h>RX��:]/�f����,W�6���h�'����i5>��fxV�r�g�tC���Ͼ�BX_-�l�[cw��� 38������w3��_�\T�]��m�O���A>"���-�1'��)����5K��g�ֺe�Q�9�z)�'���0��:X����b$)�@�
k���K �_�FV��<�f���c$ؕa��%�[����3=�< E^2���Js��1$ �4�:�,'e�w0b�r����W.S��kg���$��H�<p	[}Į�N-��@Cq0���i ����C��%���8�Y�s�9��`���jdD;f�nG%N�p�a�������}�G���rx(P��\���`"�툰��'�����0�Wi�&ɮ��H`q��`<!uN,�;F|.B��st% R7��Z"�r$�� ��z��b��-�ͥ�؃���Y���xV����ͲW����F]I���y��NtR~	��w�m�*��(�r�f�tc@��s���e��7����{D;��1�V��	; =W��Bdj��u��7_���Ѵ�xݾe�,r�O��%���R��C��w�.N��y>����A�lM9 ����	I��?%�Ha�\��U0v��6t)�o��ꭳt������h���:��p�pZh�.X�/j��'
�Eo��y��Uԅ�8�X�	l���1O�K�q�5������-��e�dr��^�;�ğj��j����hğ�6d��g����?ڗ���#����FĶW{�FÔU/�B�\j|��R��ҳ�X������]�v~ۜ�<�M �>86�A�'��=۶��rU!�$��ln���ӗ�j�w��1z�f�$S���!4��P `5�
.S�H�ǋg m�-�v�ifS�or`Q�ѓb��{j�զ |B,��4�q�[ȣ�BmL� &�h�����Sג�N�bZT��ȸ |ߩǺ���VI����6�:@չ��;�}a0�_kp:aM���(�N��Њ�s�[��5|��B�VG��m&�f:��B�5�Z�ye��hnp��fG��~�<(�a�u�I�XS���c��`#��iݷ�p~�"�?�2[��Ҧ������A`���
��Ea�XD(�l*�+��7�K~���l� X=N�xS��1��	�
�z�h�<I"Iמ����`�pLx� %��R:���>�4O��0Q�.�~�m�Ƣ��`5�K���ѱ�kXl/cH�E*�}탶&,؆z#�LI�(_*���������J횃�<�a�}i]
�iR���>[�{N,�.	B�6��)��X�_8�.�~�)d<˧G�w�p�P��/3fDݻ�2�^�P5�A"m0�v۱�\�a�C��K �:���w*U� �k�?����ڷ8�nQ%�ґ�y���=N����vLF%�<v���p��g�6�40	��$�\Y�>�ܐ?	�T`硄vl�6��c�/�4+q�-,�x� ��R�9$7����l3�z��Px�Q��˲���n���E��Y�}��mh����>��%������W[��o٬3���X��p����.�ʕYֿVe���O�7���%a��o~�e*uM�w/��:����g��hPz�)��^�>;�g&�!>1:�!��p|���3�87�@{��r͑�̟]~"��K2=��=J��Ihp�
ǌe
}�� ����52e�LS�?�AWە^�N��PzQ�L4n�����Y�j�V7��W�bO!NO�ZZ�4�r�x�3��j�]>��7�P�&�D�A;�|����p�e�f*�h�,Ӄ�P!͑��Ev¯'Q��OK��X/�,ņR��� ޜڊu28� ¸�ka ����P�(����,�:�Z~(�y��X����������
`Xù�6�6=z�B�,k�4�Y�l�ϑ�����G[&ioHp���x�R��M6��GD�>?�xwQ4��#)��>�}��-�Ef���z���j�E_  �<�G��)SvI��+�݀�k�4�!��&7l�g�O�J!
��IYg4�e�e���AТ(�m�(��X[X��FU%�]�wߍQ}^��G�xҒ�5��z=�k��m��s֖Ej�h�2��G�8�ۉ�8���68hw�ɊW!*��z�D%�p���3j�ݒXl���-��5Ӆ�����6Ӗ���{�E��\Cu:�y[V3���8v�0Y����R��=Ao2�gP��P"߯F�%!TcY�;K���c���6H� �XIAB��u�f���,���(؇��;8�����XPNZ��#�2fk.ì��6� ��U>/~�� �@tkI�ۛ�o��d��Z�0R	;���Cw�r�6k�ƨF?�p�O�6������$��&����ǁ���6�G+=�-Q���Q��Ƀ3�;G�rb���@`�'p(]��Y�^��?�]��SӜ&���5@t��/Xl&k���)� ΅"��4fM*�	.�Tx��~V�ѐ�{� gd�>�7=OYs��in��0{ClB�߰+R]xx��{	�d��T��O6�jHCa��D���NP�Ϻ�aT0�</�Z���tL�C2�G��+n����J��\u���9~�[�����s'�R�@��QK��od��~�m�����A��9�1J]W!�(&�)�Pr7, �l,����>c =� I�B@�'��T�%�}�K�W����A�VOE�&ʡJ�,^��R6�4�T0Fh���;�%�N�����đ��NN]>�\�
��c(����e�s�vm}� )�MTN��B��M����;a����@���Op6�OF�Lw�Vn����"-�̣(�eҍ +�%��e���w�����]u9�����ko��n��b(�����|�AͲ���ݓ�cQ��U+1��+6��d�s5�F}`I����b�2���&�eLS�u��r}�/Yw��D��) 4+�`�cF6q�=fYuy����L؄ެ t�x��B�EN��q��xR`���[yV9 6q�)q�bam�Ũr>���1��>9�rx���'�]5��R{�>��$Sq�����c��&4������?�La$l��z�/�p�綤-�����g=��c=h�� �4��V!s�QW�
V��tK��V�M��}�eZ��)h���C$t5�>Ң��Ε�q$\��.��t	����kuD)R�Z���@�4-�V���_Œy�� Zg�ͪ�;zfgsQ�i�k�N���p�U^D���	��͑���L���Y R����uI����v��JL#�o��y��d}���t�ׄ���p�ކ����৲m]�;>s��aG[Ƹ�o�"�>���y�
uzXh����(�� � i���2G���𡋡ͱw�����נ��S��5������f_���ͅc��+��'!����w�
�1�K ���ĝ���ʇ���8��%B�*�� �<���������L������*%�k��1��$�H#EQ+���JRz�����f�r!�g����rD_�F��O����Ad��9D�rD����5#��ǴBN�i���ZC�P�_���c�@z� �>�0�>��)��+�����u~�/JL�����)���9�|*	�.�L�7=��ꮚ\q4T���̉�4�%�p�'��2����������4�K���H��Pbn'=������l?n�~�i-��Zp�F��*�����S�`����w�.'*U�`3) r�cx%J�״߰6�(�^��>�([�':?X�Q�q������h�Q�]�_F;�2�0�W*CcF<ͱ[�)-�x^2��n�1��&��׭�i���¿4u{(2���K)U�B��sl�oվ��`�*��D3|� ��9a!�P%�[s�$�G��6������	�_Wо��2xS>����)��"
.�}��<_�@
���PCpq��J�������%Qr��t�𑀠�DK䀊�t���5ޓ��,!.�7&k�+"/`-��ɢ(G�\v��R5�� �%�"v'mod���O�x�f�����������z2�ϱ�`��q4�)+��|+x2K1�Ra�i��x%����*/Nk��|��NQ�"+��f�ߠm�b<^������.�jm�X׌Zw���h�;T��aҴ���V�ܓ�pT��[�P1�Z�Z�5��F�N�dUw�����|��cE�1ʾ���v]kPڷ�҄4�6�M��Nf}��TY���%Gg�(ް��V�$���O��C�Y(FF�P�=l����V��{���r7��Br��_��!��=��7��e��G����|����\�<�-� ��@��q�
WVY��q����#4������c��zE�=V�\L��5y�io�cM{3*���f�uXHX^��R@��:��uCM���+Gd	�K=�u;��$_���� |�|9����D� �W�U�N�VK�M�Ň���z��~C7냊�_�'�s{�:����wfE��BmE&�10��%4&�B�l3��X����������M禈�j�F�b��%+J��Ѷ(� .�-�5��#���7�g��+�������P����\�Tc�D�5+�JF�IYv�^��Ỳ,Hy��~�ʭ���q
��D�T!���v�D..g��m�E5���:XҺY�6AѦ�?����
@dL�}���e�W�¼ij`��x���eBu���4�cͼ�O3���pk���R�n�4簎��̺p���B�	L���$�)�g���l�u���]ir�W߼�T8��b�?��ťl3�\PM�W��Х`��~���O,�.�׶���m[Ԃ� �F0|�mV����M�s�����_�36�K�x���s���1�V\��7`��D��:�I�wx_*1�^/�hR-Ϸ9��쫷H��휱4�%{D-�5he�t3y�K�rcgT�:��.L��1ǹ�j�7�B� R�X��d%�v�`�tN����W�˫�9���r�blT�o��#7VS�^ڧEO������[�	#���܆�u܌J.��$�T��0���3�q�O�!(6��� *?���m:l���W��~�e�	`����`���nDJ����d�������U�`�W��Օ������e� ����w��~���#d�}���d��(S&#4�=8�	��F��p�I�xiz�VFo�)�M�[��nۊR���h0a���}5�FU�MFB��~�� ��b�Ȱ�+%:"�;��o /Z�U�-Ce��W�Ögb0���Nv��%m�+�>��-���q�;g-ªK� 'd��["��~��*]���0��.i~K�ގ�F،����L?�=ړ��>��X�ƺ+#N��������b���AȽ�|�dCh ���𯚃�NR�uu����7끯��뾜�Ely�r^+��y�����fv,�>��U�g�d2�c�h0��šMZ/�%�s�Ɩ2��5�r�y�*�b�}�L�GaS }wn��5'��l�����(S���AFn� g�l����Z��(|��]��<�ht
5���*%S��=��"hF�VLy�������_�0c�~�t:������c�1�����V� ኯם�����z׋;I�ϑ�xB��?:���A�0/(Y�fx�8_�D�-�"�$�@��j{�E�6[U�G	��%���og@�g�mc�M?<Z�P��=�Ԟ,{BS�)�t_D��YUh������k�d+8�����{�z:�A����2q��Vﬡ��].G��w���v{b��ﴝr��\�"2'�Ea��:�k�N�ÊX#fb�Ihܣ���v�־�~�&|Zb���xt\�*�6;�Q��e��"�[�ؿ��d:�;��Yn*��%!U�=h�B6�G	Jl��f�4�h>G�|N���gg��g�C�5��(v؎u�J�k�9$�M�s�Kjĝv�av z�!�˱��~�`�&�?�ui����Aj�e��@
�G[%c"BN�w�ݱ���ez�Y�բ/"�K\&��\�%������"A�z�*>۹'��ˑ���%"y�As�=8Pb^|�lI
���k�����0��C�j�����kG��� � �����l��6F�G���=|�t�g�=_/t y��A����Nu6op8K,8��>�r�Yt�6�{ȺB����T�j���v��gy�>�M"E�|�x�@�l��ܻ�#"zx^�:	B-���"Q�Jc��h=��X"� �/>,�L��"�u�d G-[
�~+�^��9��`�����f �4�X�	�N��55G����Y��H1�V���H	��b���1��M8�>_]�+a��S�{{|���EW�ҋg�N� 5]^D�N�\�!���Y_�h� m5}��W�N��r{=ʬ.��S0a�@������Q!�&'@���
^H����[���q���ء���Yv��a�ԋ����롡Y�����Jr������];U1Na�k��\-a9�l=�nm)���.V�n��Q��̧��U�V�q��}��#X���?�3����S��e E��TD����:�9v���Q��ZŬ
���!vXNU�=~D��X�K},Vo~Xi�f�܆�-w�������]-c��ƚ�a,85eh��Y6/�;J�]�Y`��7�`#�_5�l�����3�/����V��2_�QR��g���M2�HI�;����R��ב;��ŢȒ�Uޔ]��(�Kl�
���7h��W�@���Kv�$�9L%����f/3��������x�k
��1u���N�n;�w�9.]�p�>Ȣ�.��řT�{R�3@���ar�UQղ}g�ȯ_�k�x�g����<j�w�2��E��e)���i"p_HUl��Y������D�����y$�p�}��/Y#�b�y�ҵ�5X�(?���Y���ۄ�H�u������=+�N���bJ�;r"1K�p*���iN��@n��7��O���?1)�-"zN5uE�� |�7R���R���� ���N�wװ�^�T����J�Y=0Vp8��g�͡=
R�
��D��G>�$�0�s�x���J7�v��	w��Q��K�5(fh��ׄ'�������T��p	T������"Ｎ�:�AQċ�VOf�*ʲ����5�vp�|U��OE@��&Vx޷;�.�0).>�S-�.<���4�^ӥ��0@����!�y��KL�[VӘ�k�9]��BZl�D��ý�\�/��������yÕF0b�q��M�.m���2���#�II� |z��r�\/kѓ���@`�gRyߤ���G=�5���=���nT�Q
��h������Q����:�7��j:���^e��eꍻ�P��KA�퐳#���h���\V�mL���v�ؿ*�J*�)*�|H��'�š,Ζ	�څ�rr��^ì�$�i�)t�{��p�o�0�ޔ��oԸ�ҡ|_�.{PG��R���R�eZ#1a�1�������_��(j@�O��ǎ��	ي��m���W4]�O���i)��>�S�l���#��\�G��^���z�#�p�7�̷�e'x��;�u�f��K�ql���H�%w+'����|� ��/"� ٧>��}���Gp���s�FC�h�lnv���)�mmy�h�uP;�����<�Z�]lE.�3����@�$Y�to˜v��/]#��)P�]Z������l�-�b]�6\]Oy�/`���U�.vC@��w�[������ 1cT�n���|�������O�=�b�+�/d �]�Yu�S��l��adZ �O^��G��Yu^�[D�_l֪_�B;U��2��I�t�e���h�w�V$�u��挷�:�5dG^��ԯ
�˙�K��Re��5=�3&��W���ڞ8	�*N�;�3^AG�g��#,�q�;�;U��d��/�l�g��L�\ʄ ���<fE�2���z�1������W$����5_�pT�QP$<�2�U����
f�ꛢ��-'����Tk&���~��H>f[���1��b��C�w�x��3��D��=UF�
����o4g:��t�d�j��Q�sM=\�J��O�d���B�X�5�#� zT�K��<�)X��ܙ���Uo�A'G�g�����}[��3#R����d
&��cv���AN�d��Jq���_����BA��><u��t�3���)=`�[�lM�m��'�9v����X/�F�c�#��)�f9o���i=���V^��A#!K����� ��_�O�|0C~�ss<�I�޻������P�R)�D�£�I���{&B
��qn����*GT��L�9��H���Z�fr���7�H,�}��߮7�/h�Xz��*?P=�Z�^ ������PKK$���D|��Jx���b�KZ�S����|_t�	��c%gꘚ1���+���y���z��vՃ�Ir���.����^G�k�l��J8-��ܲ�G�u�{	��������܇�P{����V�����F!�*=bs���˧�7h��Ԉ�N~���Q��(ػK�4t��2?nmMC��m�/>�;sƩ�J�~ ~ӯɍ�\��G��E�M'�'��J�o��d��CS��C�g����/�<��#����R��8��*�d!��@>b�蒂���]7����?«�Z7���o�*է��Wg48B�����[9"6Z�=��i�2F��ٌ䣽��@ *���k�eI��l[k�����u���5�i��t�\7˅P��FN�_R��2ZMg��l�K@��"N��d�� �O��)w��\)����*�}C��)G�È��n�ˆf��#��K���M��l^�����Ù�I����`t�͹��C(�o(������*�\�E1��9�0 �q��O}�%l��.��Pu!4.�tf�Mq�D8�I�Ѧ� ��j����"��#v��ܦ�������?7�{���ZJ tC����)N8��dۊ�-�u)4�;�+)���q���}�΋tۿh{e���՗�����|��O�lS]&z\�Ρ�h���$�߼�pS��"r��ȥ��[ s吝ë����Cݿ�?�:�<����`u��O���Z��CR*Y�2yt�~��� <��!vvҮ�ew����*P`�-���� |�[�L�����b����R���L�����j�Ŧ��/<eSҰw�5d�נG�~}��[��[})~W#�Kd�Q���?�史|@�&,���J�Fv�m�Q,�~��$����j&�~�ªj]3��gn�/z>��+zܥ�&
`�_Gp6�S�.I<�ů5�;�Z����f�2��^ܬ�����gH�!]o��\�7r^����Y��¤�+�f���*��נ@s=��_/�Z�AF�F���"W��@x�)���*,�K�B�oe&���Q9a
���(��yT�1 䐳W^�64��^��O+�\ϮL>�v�t"�TY�_J�N���{^_P���E�[�ȳ)�^l�ĘPs�=�TG���Zi�e,�r�B����k2z���O�Ɖ/5
p$��G$����.�Ur�}n�O��#ۇ\�w=L�o-�)-N�.z�b�D�О�(����&�1vLngb�1Y���c��|W.xǆ�&VIl��P��=Xc�OF8���bѪ��s���1��Fo��d![{��*,�������<k���C`�!ҡ��]��v��Qs��.<[�,��Hh cpf̎c�3�xf/AG�Dɳ��a������<�ǝ49`0���{�dU�nxI~ը�ן��e��t���V��]��x}ǹ�+�'gN���k'�V��{��{��tB�3
�X#`ԝܧ	�T\L<n��eO_�37�7���'��� ��D��B8�Tw� "����:�}�֢������*��$)��^��;�)v����gZ�����NsjƗ�&�紿��vh����R#��)�����b� �Yeh~I�:eViF!ҭڊ��^E�I�L~��m��6|�QW�#g͟/bp�W�4��ZU�l�o{�L�Â4"KQe4 ;7ɀ��O�h��-dI�����b`;��$�)�X�wo�mw�9�1ɏ���U�����]�����p�{�R���>�`(��]��$ǡQ�MZ*yN��9�+�'�d�k�w򫂌*�LZsy��t�ω]o��g!e�l<�����G�x��\�:�1>��
x��Fղ���Ez�YԿ/��<�`]�j�M2^����N.���
��H�u&N2X�Խx`ҵE1�{`�P^ �$�T�x��߷��~��s��V�]
uO�?C�۵Io��]�wǺ������j���'9��bqo�[L�@!�]��[giaɼ����Y��mJ{�NZ+���@�U@H\=�t`����=� �L[��^���=�Li�bT^�4�ȫ����dɫR�b��B��`'�zgncm�Y��ٳ	���,�_�#�x�Ӵ\�������T"�ߧ���nm�B�dۇ?`������T��q��k�<�� d[vl�Sy�4���&9 8YB�bf{)���Y�0Cx5���}EZ�/V�3�;����}���%���D�x�f4`��e�e�����L�VX�r4�k�z��xA�����Az��/��9�>x�6�)�ܵ����@��yת���yXF��k��. lZ�F����"��X�g��"=��Kw��d��ǅK�4�j��S*��D�)���9��8L62*QG��Ey�hdQ�Y&�ު(�~�9������nʃ dͳ�N�l�k�W���\HC��N�/��T�g���,�t°fQ�/o��I<�)i�ɕXev7�[�'������$&��˸M�[��$��=]���D��g��˦�O=!�ɸ���3^� A���<.x����?q)�+۸D���B':�f����˸�^?�cb�S<َ˕�8O��t�$��$�Eh�F:^kf� ��c�y���gH�i�}q/��d�yP��S U��Ɋ�+T�h6NV)ש�h��J�+��� ���x�����U���L&�8�E!cN�U;+B� ބ���D���\^ou��Hw�������50�ol�c=oГ�1:�Ǡ�>GQ�@��^��Xl_�q1I�Y4JL��Es]j,{&���kos�X�ڒ�-xߜu�^,�Ѝ!������&��7�򹡶�J��Y�wH����T6-M�kd��2
"��"v�*�Ԟ�*�g�R�Z�M
c�֯x����Ldf����k^u@��Ф�B;����c���SO��v@�ҝ]`qw�e���e���8������bG��(%!}=��=��M]DQ)�U/~�ce�|g�¢��U9@�=�_�=��!U��E~�}2t�T�Q��1�������?�b_���<gEr���Ƞ�>��=Nݏ���zL"�rV� �`�.�q!�/xTb�I@qA����:���+_���撏���Q�h�������1m3����w��Ed6l��u�1�\�E�hP�k����� x�nq*�fN����:s6�M�vﹸ=���h?V
��f�ԙȗ�³Y~���&�|��v$\��I%�Ț ��Ň�lh?z>^�V����Q6�����N�S�
|�/"��`��9͇ToL����۶k�eP9�;��\�H�`��fZ��b��]j]ŭ�h�ܷ��=-���}����.SE4"1��
�t�r��Q���or��6�Lz�!��$�	~3%�9�55����1f�q9��+]0�3��09^�2A'N��$I�Sp����G(���P�웒'�v��q�C��x���������;i�VE�4\#�yo���S�HEE|#��aG�L�tS	�Hv��9:VX^V�ή;�}�4R�EO�F�A~�u�����+��e+RI��L��WhuA��P���L��~[��k���X���`��QxmYFz�I0[B��g�Qw��|�ڥ�Rgn��}�q7�O)-�h(�#��4���a�B��҂:f�}���q�����g�;��2a�����B='�+)�X�=8CV���r{�<Ub�)�8oQ�t�J���Ȟ,�K�z=@����t� ��J�E��R$%/Zua�d�t){tdz|U�c�w	W���Ck�S@�4��V�7���s�Y���J���%����T���r���˿d�a��k��>�8	c�7���،_3V��
�k#��w�!fDvT�[\�ivo�28ؙ�tZ�u&�ed�����t�����;�� ���d	<��2�+�9ѽ����w�
���T�e��������U,���$?��J0�?��֖
Y�+�mr�����୬P�^����$ړ0[S���A�͔�"���o��X`�j�ۧ,���� s�D5O���e���-�2�X���M�|����2�<W���9.�w��X�gLVR�b5�������b=�������zG������*<Α���"�����(<̍P�~V�P�O�z m��q(�O�g�:�վw��vY�Qx��VP_XX�k��Ԁ|n�1��?��������R��!]��!�H�`U}f���<f�V1�ݞ��[��k�C�ta+��]��,�ے9����^Ps�V.�� �bط���Z
��"���L��/f���ٟ�+���f���@���9�0��SL.a�#G�D���(����TE��R1`�������T=0�L\L�:)���T6��������� YD0�9 ��5���]:+z�����(���mO��Cȍ >����d� 1fa��*
�a�p�n� ��{��|�r�8��N�T�RڎL�;�k�F�����������c�Z�F�/��N���&�YXL���D��v��C����y�#ǲdOV�[r��۹=��o,9,�s%:�V�v �'~	�w�`���}���4v�l΋�8�#�j��te�ժO|R�����Z6�����x��hw�x�����o�Q��)X��tЈ���#���������#ͷh{@^n�u�i��f}�ZW��=�2�8��X�̣�$����$N M��V��>J33��b�]�<|@��t�+끹y��~��Z+MS-��P�H@� '1�fO�N��\�l��;P_�\b�]�!	[E�]8w�Ԣ�V�e!j}F/"�Y5��(�7ҏ
��t!�f�d���nӖ���־f<A�ӡj��ѽ� �B���%T�^ޭ A���[?��w��f*�
�u5Zrzބ㤡:�Qr��@Ͳ�-oP��	 ��7��z5�POq�
mN�e_����i��t�N�^��M�ov�$�У��URT�G�
nOYO��^?��ϰ���&��8�<����w��T(��"EyL��G���Ȟ��i�����{�v�$Jt��ȡ+=%��9A'zM!�;�K=����V�h�o��eb��H������Q-�����R�/VI�� !�W����5�z��w�\N�)��ph"� �k�il8z�<�����=�З)mLj��PY�>! X��o��}ja�h�Dv/?���`��n� r�|��t)��Y�+��	��]�s��	A��s`N�a'�_���A�7}o���V������{����&_3��
�7<�dg-V׻O�/�O�����p�c�m�n:��= �7�ᨮ���^p���mqn�:{�(0[�>))���]W��'j�:BmᯧP���!��TF�]'��=���)X�:=��"O��BI-s�����C�̡i�[9��㫭7�o�rZʁŉ����u�E����_�F�0�C&8�<<���B�-��)��q�*���7�&3x,Wn�g�z����Q��*<��_/��:0p�E�y>|
�j�.9h���3o�g�XgPF[
������ߓ��֟��v�ő�,C��}��eՏ�Z��fƱ��j@	_;݀�F�hhl���xG%6�/���ʔ�}��o�O8��}n���Y�P��cNP��t���_P��Gn`���%ϰ9�? �Q9Ar���.�l�� �B���귯3��w�hŁa�8�J���g.��)�Pđ�<G(ֶ�e��`a�Դd��}�9#�Y�B��^�5��zF�0�X��].�B�[s�Q�Qt�`�G�_�����}��Q-���"K	��W�,f�H�K�H�_*�эw�V^u�$ �A%(��D�W����L��vz�eD|�<��D�kإ�1�⇥�rq�����5l��	^\3;��	��(�)u�D�����]����]^��UB��;�3sϿt��_0��z�����-�j�$X'�����So���U�-0k����΀��?�mu��O^�g�Uqj��N��lhE�����M�5�!N�D/}�������C�z�y�	����;�E��1-��;�vb��;!���9'w�<V�:���'�<NCޢ)0Bp��g��J��`��,C-�����H�8��v����'�͔���q����� Ȏ�e����f���w�W����o��<G�'g�4�m����1*�?��M���W��0��\&q.#屿���/�c�j�.,�{�J�3D:ցR�>ث[ۯ��]s�IF��f픐��X�*ըuSp�����h���0w�_���R� _�d-Q!N&�P��?w2��_��H���F4__��pg�!�� ���~�ޖ���'�3q&=}�z��<(�2��]��FD���ޯjګGJ$�����5�էH� ���]�}*��"��VoriEۥ%��M�]�CQ��4Źͳz� ��;W�<�.b��p��4K?��-����i�s������O�[Q�.i[1gF�W���r1wE���n9w8_�bF�=1���ǈ�ϹL���Z'qP�:-��(�ߦQ���@������%:�B��*��x��]��Q�T�\h0
x4τ}0R(�l���K~�P�Rul�����7���#�S�	}~�Ϸ/�q(��0����6�|�K��o]iIw�c �s<?��PJyt���d�_���dn]��T����#����,ma���� ��ι#D/p��Z�W��ue�-��9�3��QY��Jv| �5��U��RD^�0�w^}����r$t�;�pd�q̲Zk�w����@+���1R��4'�{�y\��cwV�	��kr�B:�xo�@`߯�O�T�gy��`ׂc�18��Y� \g� 2�Ep�FM
$��)�$�Z��'~��j��+�Fzkdrl��2�6�����Y�j�TK�� h����>��sAo�����=����팆��|W�&�z�F��{p�,E�@�1���ԥHw:؃�����ʠ�$̩=� ���Ќ����Z��)��ڰ3'�Gw@����be�3�p�F6��=$��f��ߤ@a�K��^�� D��أ�ڙa�zw<����.�(_e�l$j��0�9x��7j���	{9�Y�gOC�D/�Y������0�ˁ��iD������ϼ[/I���#fNу��a�^�}�i��~��h�z��<Z�O��ŋp�� ��(O�譭$tw�M2��b��밶#߳�N`�SR�H��O;�x�&������N%r )��i��������D4��j:�ysv��e
�_�+��̙�2�>��4<MM�hw�u}���gC#�f�Ό#��|V�S���-��%�����~�Y����{Z�B�\���i۔n	ى-���<�-�5 j��$q���� !$Nt=�|�e�	�[�%�;�Bf��r�����h�����c�+�����
	��c��:��A.l.X�����?�%�ٓv�m����~�aZ���P���v�9�^�38�F��"�I8��--�#����im�mD��6ia>*�b� ~<MK�g]���tO��aI��cS�|�"P����o^XXH�5�H�v���^�輺��
G����Z��|ۃ�,�j=/���dԕG��HJ��]դWO]i�Y�`j6?��?NīIt
#$�*���&A!���������L�3>�]5Yn�C����p;�l2)G0�������K���?��7M�{0��!�_���ң
����X��^D��=?,@���j�����~�6�~D�c����3lkXH����|�޳;֩�qȱ�<Iި��vm��U��&��)��)��RL�����ZZ�e:̖K��'6TV��2P!h��cY���j�^}�:>ǃ��5�69$��r�n��G�:���j;�F��Z�H��wj�wZ6$5�juG�F�Ʌ�����c>M��n�:j��kpz� � A�y��� ��ay?�:����Q��͟5�
E��S	�:�l�|�=�0b0.e\%��^��f��[�4��mZN��Z�AZĈN�僿��E�lmϯ�cQ3�
��V��m��+C���g�H��G�7�7VٖQ�2"���;����}O�P�w�ܦ�Ah�����w[p8��O)���&(�j�ó��>|Z�S�7���N��:�������F��`�j��U�b���7���m����Fj���1Ɛ��l�c�+	M��KR��*-��F�/h ��6i���~�ǤV� ��S]��P�PGs9���$�}DPB"� H�D�q��_"Шu�H+ݍy2	�I:�T���$y�ć�{��6<{fZ%٨8\�r��FP�զ�����u�A��&�U}���*@8�l7���N��.:��~`��n�Y�Sۣ]h�@~K�����FZ��E�m����, J�:(J�2����e9%����CnҞzb-ۭ��m�T�F/St�l�e�iC �w#D�F�������g5��rTt�Q^��I�d"��c�7˧�.�1	�,���;= ����K,~p��X>��^�
�C���6�kƮ������"�q�� �8�'�	�c	�U<V$��͘W��)�����n�[�� ��W�X9���}"��լ_@Y�����*~��
�)?�ɇ��٤ݚG�`+��CfL�0���J�y%| ��e���ݢk֯(3����q�=�C��f�y��U^a�
�F�6~�� ͬ���?��-r���v1�)����l%ir��,���%���E"�iP�Q���ޡ{�����P�ס�#W��!����d���I(����8����齆״
F|���мu�6�F��s��g<�	��MJe}&y���4g�K;����G��0~�9:=D��PѠ��@�b9��8��
��#O���������xRO(���9��N�\��I�:��n�D�xh��X5�lC��.YztX<210���f���{碝����<G2p�,���ngGq;`���T�
��쉵 ��'&̺s�j.��	
z��h������)з�t�G��`5j:����	�@����g�3mž�_/�>��U� ���2Wt�<�8�ZMTL6'Zl3YYG�Ι�����}����`̐"���S��$��9�gV;1�t>��Y9N�'w�w�Z��R�I�����\�EP|n}4�+"J��QA��2Q�b�|[�[)|�ӉYS�L���?eaؚ�u<��Af�	����U�� ����-ډ9�󔝴��m�X1�]K�;�d2g���E(�T��;�C�2{ֳ������
�F�T�fF��b	m:I]�H���5ө�@��\�^�2s��hBĪ�rHG����i�ޕ����[ߎq~˾K�F�Xq����zs��@Zn�瑪r��ySy�7^�W��1i?XQT��Fֈ#�J�ϙ�B��Ś� a��^O�&������1�h$�z��ks�zc����,&��fe&2s�Z�Y3�8�q4���x�r�p��&|������DZ2��Kx�5�F�,s��vr��|���r���3K��I�!),@w㳯e�&-�1xV����J�1m�B�1� ���<�S�¡���)�%�55m1I����9l�8� v�' �7�=!Rٻ��yɅ̣ti�`+J��+���<�Y��mG�5���1
V.HB)<˚� [�0K�բ�����_�R�dm�#�˾"��`(cCcg��eԞ�ٯ+S��ed}�b;4�z�Ӥ�����$)�=�֠�/dwU$dcI$}<
/�i	����EN{΁����6Gt�6B��j�M��e�A�T��������d���+���ۖ ��������8�����i,�_��66l�`��485�����Ղ���n�m����&�`4�
	m��m��L>{�Y����`�a�`�x+xv<��P�(�}Mo�͟l#��;��sï�VE�ћ���.���4�,�*�,[�Zoq[��Xn�������G_��z�a�*�3�WO-hI�� �T��o3�s�D
���3��4��v�"��F���8�C��G 4��
���Q �m��`_@a���l�}ҩ�my�r���?�h�=>g�J�s)��
=�Q�$��ƭ���A��kH�\��Ե�y�f�f
�����M՛��aQN3:\���@�8�̩:wEq��p�������g����k]M��	�=�����u���
�T9�Gr�Ҝ����0�_@D���`O�;ʈ+�$��ũ��+��f1�7�P0��X������rY�?�`� �!$YJ3#�~����2a�Ѽ�N�(;��P<�����69k�a���.��l��M���$�k��0�6�Q��E�$�n�j�\#�/mS
�A�g3�$$�0�E�*�%8vO���<\�,^%�ձ�:���8<�n�.���Y�)8$�Vu��"E��rM�N7��0'
P�΅�Eڅ/�ryИ,'lb��Em��5=dI)�}Ւ����[�no��3ֿ�{�����V�W:�0���~h-�=�'�?�:���ۿ�6���W�Cy�]\޴p�ɘ��`�\�e�IuԶ#�K�Ls9������WB��~K[�(g�K�+h�$J�L��O��2/�	�e�p��͌����EԀ9ۼ���|�8M���%	-� ̄֙���@��.h/nw*��'巘ވ(?��v�Q[hqa�F�Q�:@)�c���D�V��ETo�LuKV-]HRԶ	��.vRG����X�Za��I��Aw�t����9a�7p���<y'X���_���cUך40�0�*p;-������������_�5����y�I�v��y�V)�c�G�ș5(�������jgn�g�(��ao��r5�aW^��Nǭ
Fs�A��y����r�������� �v��T(U�@liU�T��Į�!�#a�+�������i�}��(y�}��7Y��n?F����y&1'qc��v�*p�I!����1۬�|�f؅�*�DL4��7�s�A�8ȅL�c�ɧ!���+�.��]4|Cź�|����@��o�T;�o;0J�I�W���l�
��'�=$�A0²��8sY�$�^%�Yc�Z����cޗH[�+i�AuGP�IUčC X�F� �_�?�9��R�ә�Nu�����b���mS�dG�h{)���F3�|hT�Vʏ8,���V���JoL��~$k�	m�
�cP��O�dW�4\�A8�3$2&�^�d��G��'mY�`�1���G��n��j�����m�sY��O/��e��b;"G^G��C+��V����^Sj����e�z��c��S˒�:)'xo�N�?�х���H��0�/��%�1;����S��>w%׶{�"[8M��p�O�M�d��,^��!}G����ld<>f�u��G2\�>�W�i[����ܓ7\+�m��C�ߗCȨ/�~�K[  N��{L��^����C�sӟf#1��$k��O�J#�����{�7�۹R�i}���:۵PW�vYϦ0h�����h?.\FN=2�-��	�����a?d*��nҠ��"�0��#ͫ��8i�ZH7Nׁoޅ���l�����,��*�S5�}��
dS�����1�J���� >b6ƁG��#�m3F���?Y��]6%#y���A	�adL�pnT��^�x�s�M���q��$�.�[�虳K�p�����E]�x�袛�VL�
Z� ���?$�6<e���]�8lx��e}?��U;u���O��6�{��5��}BS����n���(Y[f���e�Dzv)̠�~�W��co�zr'�}RH�'��$���9�P�u��'�=/���{�g��f��fg�R�iN��d`��gy�3`i[����Dg����ᣁ���VЃ�={�h�V9GP�){�}=O�X����蓗W�l��f-���ZNH��=��&:�˕�U��9���ex�W����/�,��[��@|�~0��9�Ŝ�rH�2��rq�#�˔�SD����k�j����gSٴ:�<!���9Z�k�l��ТM�H�[�$O��|��Ʀs0K�Hd���2ws�
T}.T)��D���6�P{�Mx1�Έ�#T�8�����t���� �0�q%fšl�
�`2��D���E�
=�դxe��-bN���X�j|p���[���>!����bT��+�^��n�U�&M��X���v#~�����ڀ��DL�~ш�ٓ�@w��A��TUSq��$i�d�n��>�z�,;�Q�S2mə��w��u�<.�������8C����6����_ �>��8+ �q�3$> �~�D�Ƙ���Ih.UEEx�'�^�H���q�e��n9/#�W��q�*ۣ���+�t��X��9�� �m��0�5�֯<,��w����H;�nq�rTT���b�~h���aQ�c�V٣�YM �*�da��� ���E��������Yd^�ƌ��E�/�:4�-��;�ߐ|U�N�t����_#���K���&P�H�%1���B~b�nVhy�+�Xe^��Nޣ�:�R�O�--{��d�_;���޽�e��(6�^`ؚ156 =��V˼(��W��Ln�x�����!�[�h�t?���]=��$�"���U�D��,0t��k���=dA��F���-)Zb�<�7�l��V�E/TH�A��f���)���My8g��� �:uU�I5 k�s��]�3�~�H�R��k��q������n�k,� 5r�p{��k��濬Ơa͓�d獡�6š.](>��hmB�e3<>;�|.i�>h�$��J�vpi�_��j��U�s	fԐ��pqM2�O�چ�l%�ܲ^�Dsk������*�u4;���fi@�*�X�K�'ﾶ�a뎞i����?�&;�?	�H�>ښ_ʁv����ɋW��g�������������)��0�EɁL��6��§^O�c���&[�ЌE��.�������Qo����岳�	�^ʈ�j!�˷l�zr[�E�s*�lJ��x;N���2����>6��!g�����|h��oD��`3�C��9ΈgFyō�n��1B|��,Jl��o6�\��Z��=�G`\���YE��F��{�P�Bd���f��di�2ğ��BZ��Y�f3eV��a�ylXQs���	/Y��`�3H+M�>�2���h[c%�<Q#�#�N�{����o�kP�hJ:}`6;b�����z|�ƺ�&�lE�0��ǟ���@�U"�
��xO]ń�eK�ƧmZ����ц�lo"��"�!aK���	x��x�/3g� t�osΣ�9~�x��R���`*s�
�
����$ϑ��>8�+G�/<��Zs' 2����U��K�W	y�Bꅱ�I:u�C;t���
���KcKl �m�lM��J`�I��^�MU�x�^�~n�g� �=D7��
���2'����#=ȸ���б���D����,M?�Or	�ۭ�zU�I�,50|��|�������p�c^�+�tT���������>���m*�����,��K�_{�[&!<�0^����S�*y�8�8B(2���Х8����iYу-UM����1��#ѽl
M�x��,�-!��l�t~b���:�c���d��(���}�+o������)Ւn�I��`�6r~%*K3����RM1>@<��p�	\$D�#d�P��<��BJ�,6;��<~n!�_J��~��%ǎ�㴸�@�5�ur��=�Vo�A�j/��M���2��$�.�c������Gd����gвy4f�X�}��ٙn���D���DG���<��[Sj*��z]?�KY&�Y�x��#�lЛ��"Z9�;3M���s|m��1����8����w?7��m@���nd!�A��^k����JߵG�(M-2�L�#v��:G}��Q����AE���?Ґ��ni[��'%Wm�gh3!�D�H=�3�mJ����y�':+랡�o=�k I�e�V�@G��8Q�uj�c1���k��Z]e	�� '�}9��������8�8�(��[�١�p��t-���L��2+�[?�++�n�[^y';�.��D=��	R���OUf�4*h�˪��-|���\w+D�\=�l˼e��i��s�O��6pe�� x��͈��Q���]������ Ֆ��d����+���/�0c6��I�b/^�^����� ��x"�3�q+��-w���D�PA*���K�Κ�C��zl_�h0�S��dW��4\��(���e12�T&=��i�ڬ��)Z�M�_���o�y�C˸���	;�QY�D��ǭ	ճ�IWE�w4������-!0f*�;�H� �=�A �
�x�o�1IcN.�-n�'��)V;��Ͷ~O��&a�ޯ�\�tU�3�0�Ag=7
�@F:g��(�:+�����R�7�V�` ��<CC�K&[�.�9�r>����0�cU�HwD~2s,�^�^��~�4V��¾��В
�
��3�֘hu-������v�b�����K��>a�]>��4���*�Cu�k�K�u5�A�A�̚��1�9,zN�:������A�!�{� � ���c���(��}q	>���r����7ΧL4��VH�ť�+�O���=�(k��`�J����:{��J^䘗/�~n48c�A�A�݃a�u�Ͽ��+��"-C`j���h�uг5{����i�4�7T����Uo�K2�t�QV��}��0��O�s�V��S�rܘ�3���ͼ+�+�fE[;�^Z��>���UJJr��Ҡ-?�8�5��G�06�ҟt+Q����9��7x켥��Z9�|�{���(I���^.����T���A�UxS9�XD��~{�p����5kH��)�����p��髗bF�m��^?]L ��?�B���	��cv�0Li�c��"P�W�����	�Y��c��?�K���18�V�.������z���e�v-:h���g,%��ҋ�q΋�&��V`�����~�n]�*�aWe5zt��l|]����s�&��UkYys����ȧ_�_��P٦)>u��O�\������W׎S�ɣ�m�Z�{/�wl e�#.�����,�����Z!umZxV�]��S_�`����������TP����#��Ϗ��Zj�۴{G��@�����5�ܝg��g�=������/�t���)M���Qc`���e!��.p�9��]śQj��2ɥn���ϧ2�m�r��2vAg�����1� u��:h�Bp4���� ��dpn�<�}��^<!DHi�4m�����|b�W3F�T
�t��'��lHqV!>��F��l��c@��?[?����|r��/�*}�%�ţ=iĲ�଄����6el�k&���������[�����޿�2t����x\���_%!=l���̊OP� �b(<U܂��j{�b��㩲EPI�D�s���G��;����_���x'Yd�A0K��X��dNr�wj]NX��{��З=<[��p�Nn�m�2�l&�_&�)���U�CH��e@���y/u�n�{?���$D��F�T�D�.�)��љ������@�cw�&j��))&�􌘙l���4��^�@��{H��~�����7%�H��&�4��u�kl-��HR�uʛ���(�F\�f�D����/M�Q2g�m���	5�������<�X6�� ��j��'p�wJ��\M�|�d���X�)U k '�����fL�x���>D�P��`�C���S�y�MA$)U����"��F�:˳򦽛-HՍ'<+��<\�*�"�N�?
-J�:cI-'mW�r/q�?����*��웼alT��+p�!G��H�bXT^Jw|R�qc�,m�Z��]B�Bφ-u�j�o8�-�ˬd�i�!ߙ$�z�&�TܹrRm�4�����?�������S�����(��x��<�Kk&n9�)Q\�|���,�Uwk`xo�=@�ѣ>3�u��}���Ҡ���d�Ɣ�~*��r������y���T=�z&�R�.D�>qn?�gc�3�v��]֕7�Qn�ǉfӒ��9�HΛ�(�-��3uk�0L�v('Z��B�ݬ6V��\G�!��ca����E�;����ݔt��I�� w�����"��3OZ7�����̆�٘��+=�%{�E=������IG�Гdx���t����kg�`(c���
z��N5��+�̱��F����;ŴVJj��L���kPI�A�).g��ܲR���Q$`�t35��/��,0�|w��q��ɖh��A:f����D�V	���@]�_�=�	Oyd�eDom��$V_S�p����@f��2i�gT���K-]h�8�T���`�2�[*T��c=~������J�,�5n�3q�K������h�a�-��\B �,��r!��؋���%�l7K�eV�#�9hXb��J��d�Vn�yJZ�vt�;~�U6	X} z�V7A&:�cl�s�N�ՠ�1l �	���I���lz,J����}$(S�ۗd� �f�=`�A6���V�S�D���,����%�!�SJ[E�g�Q��(�9���i�M�6ϗ�?����M.�5<���>��A���b��0L�0	A�T��{�eR���W��9?Y��<3�.�^�ߟ���SH-�v?V�Q���Ԯ�k7F��o���,�F-%x�C�/����h��c�"�!|��Q�⸼1����I�0�E)C1�VT���g�p�}��u�1��g�=�3��?t�G7�m�g1��sC[��_��.b���y��4;pQʿ��y_�P��ou�5�-,T�0�'9u� ��<��?��#�
��Q\����&�Ȱ�v�yC�9���� D��	��e������������&)%�<rf��Z��9?ji�)�Rֹ#�%�D���S����F�	�y=|��HɌ�WAbQ(V�Eh�+��5-4U�5�j���y�x\���"��2=���/:�@!h�ȱˏ��l� � D�C8G3�r�x�>�hN���D�$s~l}����jk�B0Ùr�VG̩��`�����s=�lF�U�2�!�d9oy�X ܮo���G���S㚵<�N��_|�<������Xi�Ʒ`�0~�	�:��Ov�������M ��%���W)U5���a3��-J�X٫rt�Z䜚�h�$T����`VG�O<|P\�qo�r��,=ώ��Gǯ����t��Ə�EYq�l�x�vp<��$wqK[�&�� M� �'�ݴt�(?t�PӒy�L9�j.+���ť�"�(#���3<Q;�皋��6�i ���&'X<������(*����]V�`�����5 �t���?/��8aG�7g��:�������#���@102&|CI�Jx��?��$\R]��.�[��2X�=�N�o;&?��g"s'e����2 zEf��x#�I ��XV����_��������shV�">˟y7'���-�#^�@�L	>�U}\!HJ�F��?�%��u���N�D�(�M>��GkRmNS�83�!����UV[���������D��M�r/�Y��Rĸ�[��-���[iv��k�#�2�8y��Gz�,���W:т��|�$��f1
�^kl�XX �X��Fx�P�J�����$B�%l"
���Q��{E{�#����U���=Il�`}~]��E:�+���ڱ����R��x'��b��FV��W�\��;���jS��Zj�e�e='���<I�I�
�D6���[]�K�5��	.>\}�LQ�VKu���ݠ
�3X���#�=��%��[� v$�~�Cڡ��T*^��6�"{>p��N���~|"�A4��r�	S5�k�� O�֕ƅD��A��{���x����f����cݠy=�vwmM���#}b�c@�D~��.҂�q�: D��#D���A���3�ժ��=1��v�Bx�ZxƎ�����r���5'�����FʱЛ-i<�<���'U4��m���O~�q֬��bfQejQXT�R�`�h`٨m�������5�^({��4	� �����B��K��:��BŒ�G	����&
�Ñ�>)��YՊ?W�vk��f\�O����5�T��&�7�NKo�����0�9EX�{��ƥ�"C2@�R��Yn7Ԁ���.%�%�x�Yxrs�Ù�g��,��^�'��9'���Zc�;<2I�;t�l�ہ%u��#��ʁzP��S�9uN=S��|�H"��=YK���E>M��hI eD�%b����"�S|��`p_Q��6����JE�+g<��b���{���m��^�j��	A����+bK��Ƞ�j^��
��G��l�uHבt������6vq}OW��gF~̄۲�c	�.ܯJ�vG(r���iv���#\���d�g���t�3�8�����esc!�{.?�G�z�������Ψ}���6pƪ+�����ְv��?Ev���ަ58[���[B��K�L�z�jb�1)�,�Y�I�n����^eB��=T�z������K�����3�c��Po�q`iR�$��ƐW�ΰ�,��v$���/�^�p�k�2=0C�}�	���17�_�goiXX~���C֍����8^;���m�鰪�m���1�b��偉�E.lxG�t�
gѵ���GX�<F�@f�1[�\U-�`6Jd�b��\�ME/ycWV"��C�k���_n�K	|I���.O�jZk2�u��;f���B5[�Y0�!4�z`c�s"u�q�Jyʞj�^gC$�-�"����xj��qb�v	�?��W�؍5�ۦ,D�",:�}ڇ\rU�6�e��[�%R�b�ˇ5w|�D�k��:;Ij�9�Xt,�TH`l���[�~�!ak�(�7<�|ӷ���qK�J���V ��(Yna�YE(j���{Hj��[] �0�M��rqo6����6��f�O~�������P@���R�6�@�����$�] �oO�&��o���s��t�}ضY�_�u����*
��4���`��nە���t=�d�%��AKc�B¼�1��ς�=���l�E7�`�����-v��u��^(�b�P�3��TC	ŭ_��rV��cN,G��20�����s�]��Q�$Q�OJ�~��'OɑN���*J
��2���cF�C,o#�A^Uڙ*x8��Å�6@S�1���|DO��1ņ(N���N�o�ہ��jTQ��?����I��������4&�J�Z/w���<�~D���=�t�����0�}vŎ6޴C�[�3���Y�e��0�O$�ۡ�X���r�&Wf�"�H�|f2J��]�e<1"'�,���г����~�Ҕ��a T$���,T#0��RfW�rB���>o�к�8)�����>(����>�;c*��������a͜��㏴��	�:r�D7�-&v���O�@d�����{�pO��y���T�q��9���\#�n���m�l�� ��-�lh�4�S�ť.�;�W�S��f�ぅWt��ʅZR���1A9ww;�l�x))B"��,㢻�결a���^>�����[w櫣GUW*���$ C�L8��DIk�{�*�K
�I�%�M
F���@���
��x�Z�H��Û�ޜ���ZI�,���[�D����nH`��\vm��k0z���i�-����O�R\�3�	bN��8>����x��|��H������f@%���9�賔��/�μ�V�}���Ӧf�z�0�C�Um�{a6������My�&Y��y���^^�$����c֙'�P'ϗ��j�z�-1����|�Tt?��Nz��q�_<P 9��9d���� i�>�nZ��/�;�J�c���T�wS �~���G��C�9{�C��a�k���ߐ�[�l*� |t��@x��i�+�6�:Ig(p������锈^�M�*��8���Y��k*�S��4ЬY[Q4$�GB�4�� [���|�#�>������N�QoFxX�Y ��.��FO�P;[i�B'RE��+G��2���y.<�n�_��ʒ톢C\9�u��t�mӠ�Z1&4�sF=}����f��\e�ϸ?H̲��;�r���QԬ�Q�߉!	��V��ث�g5^���w���aV'q�UKtiEP���סA����"nL�ܿPJd����P�*l�M����b��]T�w0P��I���cR��:�@H�n��l-]�$�>���~G��Z;Pj5n�Qԃ��I���Q��ϭ�	�r��1-���NIf�6��i���͢�ݵ��6[v�w�Y;����ӌ�#5�>�}mr�D��&�l!ú-\�:�U��z��ŧv�=<Y��e�ɉ����������Ihn���>:q�]��j��!?��'���慺�^��t&��då�p��|0x(9�kn`��kh'�b���r�Ȩ7�ZRf�n��A�ȕ��1e�����.��W�m���T [�tFJ�^��H�����ë/x��"J�WŽ��,a!IS�U.4)1�K����[���5�c��c���F�X���]e��{�<:C�5a7%"��bϙ	pa�ӕS6�34�.�������5�-l�V�3[��݈y��uGI�<K%/��$�P�E�R�z�LX��ӵ�z�X��.L�7����k��4-�5B8Il&��ET�B��,I(�]SɹT=���Y�*���b}Iľ����s/�ӱ=��؃��}ŋ��oR��7�[�r�^#�YLq0I��2�GD�@s�}�)��'�o����!����*����|�,]��;�;Ɯ�Qn���c�f�?Sefϖ]`�$x�� -�ʣ�>��5�짢"�\z.�3k��T��"�����!�`���h'����a?�g���F)ྔu$z��=��ơ�û���炊�K��	�P�q>aP4tH�}Z�����&Qc�G�sXy�Ȝ�q�<�)e��E(z��ʎ#v�=c���v�١�-u��(S<ި#m�(����>��tѬ?�|`��$X����lW�ga#��=��Z�m��U����z�e�X��NHK�+�����B!ڮLT^j�ؔ�B��z�A��Q�Ѭdz	ڋG���c�j������l�:J^���Ю�lyp�=g��V9�Z�/0-�C�#V���`�
��^��u�������?�B]f�h_Q�}���,"���?���}ꓑE��9Z�+�:ޠ���Ɵn�~d�S���&��2���!�o�	�gf_�y�!�WcB0p#i�L�=]�O�i��[T$���4��΢�K�Ǚ��w�?�n�����߅~P�^G9s�/ɗ	��{k�F.�@����z�iUv�Vɉ;�t�����\���6X)��^�u0�F�K�C2I��l�.����}��P������\'�w0O��Nv͞��,�Il���E�_j�b5���]�P5(�)t?'(U}.����  �,�i�����	ǹU�V��
1o>���%�ƻeF�H��O��6��[�Cj���i"?S�����hD��rU����#d��$Vj ����d⬳%P�6.��F�x
v0��r0"~g���f��G��4�4k����W/|m���=$+�L�s�QV�HI�+ǳt��+PQ�c`�M�đ�y�d	h���T1��J]�Nwٕ��l�J���2�d����ۓ�JQ~�`����,/�w)��Zb�kWJS0:�Q��W�;V�VT��F�~Lr���6���%�0iz��u�g��+n�_�[�����P@��@��t�aU�/Z��c�[�7��Rm�'Kw���A����������ɻ�e.A�<w��
s���C�lJ<���NF~��W�"~�R���E ���49���m:��$�L��,�Zo����>dwb8t���J�X�UTJ�=�>��Ro<��M��z��~��?Ӯm�ݲ�&�ᲵhwH�gA�Ɓ,S��~� �X��B���.����z#����V���������>�L�Q��f�1Jr
\e��<#��D���u~ʇ;�N�0�q]�����3}@	ntX�Xo�����	��㆘O;�YX9Y�/P����aU[�����\D�Ϥ ��01Z �@�g��O},-���j�ե�蟸������DQ��R��z�k`?��f���#5��$�'�[����&���S�/@�3��u��m�M��́@�gi0$�{l8a֥_M�9.:�5�E.�;�+E�XAd�0$F�o��m��Yz�~!>sp����̋��>��>G�.u����p�`eh�B�r�$��H�j:JԸ���b��u �Ͻ,e ���g;�`{��'����q���Z(��'��>�~����e-7��}]�II�O�����v�G�HǢĕ�SRh�=S��dS2۫�.���e�Pj&�J1�.j�/��1�Q��E\�[��x�Ȗ<�	̵H]u�%sAZ�p��G�0Iۄʒ�Vi33��]X@Fv���wa�۫*��͂8esƞ�����H�%�4�C��̅���X���pwү��bt����S~�ˎ`ɳQ��$	��	'�@]�n�%۸nƉ9p�*�C��W�\�d���z����?GB"��6������eנ_���hЌI3vP��Ec�n=q��p��r��`^C��B[�}ZLW��6{F���~��k���A����ے�~��(s��J��m��)ۭ螫.#��+ԧ.�ٶ�x�NS���Z��/X��9o]GP)L��X<���tU��dF�@5ĩ��hj��o9_�=$�6*�N��Z��+`L��Ց�iW���{�-d��0��5aC��� ��D�=�<����j�(.�����7�����P��`���&<㘨�!�x�_8�༺Gs�ղ��H�u��G&,e��.��0n�NУ!Z��D��<\f�	j���qP]0ݽ�4nvd|�݄ZxhN�s������(�r��y�*\���9�J-�[��}^��I�jj�Vm	'Y���Y���!��uw��C=I4�M���j�A��7No�~�_)��/<ÿ{`�Y������L����h3Q���JRZh�'Z.6��]���D[ #�ME@=Q7��p�std��]����j\�ë���ɲ��6tr��_����?Z�]h��:��C�Y��.^�8D��KRf�V\�d�L��mK�Uq���ז�aʹv�naٮ�'[LI�0$4�X�(�������M����F�8u��s��>%�����(1��$�T.����E����T�4gv�����_<�brM_����ƴ10�S�Ӟ��Pb
�^
�{��T'st�^�{�5�F�j,:���u���ӟ�G�+�	�hYPD�3��뚦�JX.3< Ij쿞c�Ց~eA�:�C� ���X�F�5ڐ��	x�d��!���LA���p�\O1�4�~|���hB���B@D�c�=g\R|g(�Y@��W����(�!���__<�;#s�"`�i�$BE��H��vy��e{�h���3$����H��N���[@�ͣޙg7Xx-R���T�3���Z�e����<W�6�l���埆��h%��~�V^�T����8��� ����=K�����WC��󄌆`_�~i6!�+5L��k]�&�(Ҷy�d��~&�Y��j��NQ/�>�"��.;E���XG��Xo,G�< ��-��'��Ӫ��5����X棃
���J*�0�irT�D���=����V=���ys;�t)pHt��}�3�C1�i�qWyexVȅ����*@�����:.�,f\|�E�oEU~��/��&�.?�Ę�P�%"��r�?�D��}Rf+��=R�v77o�u�Yc�퉵����HH爷�4?����{�Gm��CosL)�����	��2.�̷��@p#݊A�.��a�^ϱMRz"�3 C�?�aK�S5=��kUt�s�%W7W�ه��mB��00=�V��V�j]n+���9P�p<4�%�����P�ˉ��YW�L� 0�pI����b�"4�R���xUvX_l�9��W���B8>9����l�c. u=#�m(�$�. ל:���k�Y&��j��+_�/%��%��m
9�}郠~��I�������>��nVK���NR�F�@H��$�x���I��*��GB��1NR)�47�~k���R��c�p�<�V�1�n�R���U�RD=ID�&�w+�y���a���D�q�(1�5h�>�H�֡�Ц��
Ude�g��CXB!U6l�wyz�u����@����u������^��j����U1�dTzo�羑z��K�7��X|����Z]3x$Ƣ�E�e1������&��	��3F#Fc���m?.��� Y�1��J]��\#{ˌ]�@2�K�g��L��e�E&YŽ��	T�����~�,.���L^��/,�FB��w���C�肶��W�w!xS���,��������]�e�(��N"�o^]���/�|�7۳��xvżۇ,A�טEf�u�j1��ԚѫV1:�$�|TI���4P�߸K�h�XJK�Z�b?�g���03�M�n��̺p6�N�x�P�L�9<��,�����{y�v�u�b��|���G�'<)���/�xE�$H������;ߵ�A'S��1�{mM�i�+LJ�%7�ky��.�yj�=��ܛ�}'�F$�N�B|_��,ѯ��!]/lġ{��Z}Hȩ���t~R�������MIa���A�����O��U$�)I��)ɝQ�Yc�3�"G��w$DFl��C�/�E��'���� �#+o�i,�-�4q��E-{�kNLp�O���G�1aI�!�k#���j�ӌ�[���n�'�, _���,gGxc���'��I-�����q�Q��	�bMǿ���rL��:�=�������'��O��!����6)nO���G x��G�G0�n9��
. ���U�_&�da&�P�z ��t� �n*��?�%�9y�E�N&��lE�P���1a�
Ue��XH'JK]8�F�ʡ��9M#q n�,o�����\�ّ��I�b�ϕ�?:���h�i��9��z�;��Vv���<&����B��{@Gm��ߘ>��%F��hRF) E�+F=aEƈ��?Ǎ��'����Ae��&|6 ��^�p����/��DW����ktQQ�P���-��)Z��/1�J9>�����:���FT��V,��}c�s����k,��������Go]$�{&ξB{*�u��դ.�g8���!*o��nLc��~���_0Aad`�;���ݤ1��LVV��i���6�-�W�I�{3L��՚Z����d��<Nu�B+���<�9�+�Ŕ8�c�d	L�<�a�#�}I����x��Y3R�-�U�?�"fޜ����!C]JPj�m�H��2^�T�)�
W�-(��z-0��R��8�'y�H�m��NEuD��=W���yL7��m�l&���Uh�	�i*,P�cR�Ā���L�xH��Ǵ�W1rY�Ǐ� E�c ۷�����{p��;B�����G �h���Zv���dIe+�\4��~�����3 �R��-Y�I/M�SL*�_��%�q�_�&ԋ`���>����ֈ$�cV���S��oN���0ǘY��k%c����"�eσ�j���PH�90+�W��Ȼ���l�O���i�v+v�/V���7��c����b>�B���y���������X�~�vʇ4q)I�^2
:��x� �#��Ԯ�-�b��Y]F��6�LKL�|T����k�Q@攚c{;w��{:�Bt��1y^��q*�T���=~`],�ɝz���LZ9���?��J�[����ɛ-���H� 妳�&f �T�t��`�'�X��zk�_z�;�^<��Y�!��V	�A{@�Mi"˻n���#�����8�*(�Ø�_Sx>5\gUEB��S�i�[=�wj��}���4��[
�(B:�|W��o@���D���.C ���Aň���?��������I���(�_K_q��؎�`��|����M��x�X��r�#�C3ӾקRrr��'�\�)q�Q\za��OWB�Q_�gz������4S96����*������LI�F��q���ߡ���~�Y�R��Bf�׆� ��]_���, �"7R�B��\�W����dx3�$14zǦ�4�\C|�D��L9��qi��9Y��S�D��Σ�0^wj()K߻��$�[�ă�^qq�:t)>a�a�׳�0b����yN�5Cش�-��:���� �b�5<�	���IS�al�!pT> ��D$�m�³��#����r^F�,4ǖ%�6��� � �j4���e��3`��^/��t��\���0�햻��P�<�� !��~�psJ�7�>��q�����"K5��P���@��t���il6O?{
]���.�h�u�0ض!�o��i�T��'cv���y�M}�ިfv	7�A��yȪb���ʡ��w}p��2�\{�FA�=�Ϋ �ף>$�r&U<a��6fA��-C���j�E�CG�k\{�ꦉ6��D����㥎ɾ��vH	�>�W�l����a��X$��,$Դ_I1��k#AQ3�Z=I���#.;]6�t����zn_t��u�yXI�T�l���|P|gOa}
�8�����>�)Q�/`���a�����?`%=�u(N�&�H����;��kR�h	��a�(���'=}�/�:i�el'!��C�k^�����+�(5?�\B��x�z<>T<��^C��	�^t���Pr�|܅������x>�Dy��� ������+,At�酱V�u#�k��J�\�:r2u@��H�J^�+��p[��#"=%V��Dn��ә����v�XP�t;�}�ҭ�^LE0��d2�3�gUH]�^�ߴb�b��ҙ@ٳ���ƜE����3�TM��2�Ƕ��n��shy�Ǖ�i�⶷��΢.�0����Hx�6I=snX�p��}ɼm�]�l�=�V�cO 0���0����J��*���x��X�0�%ɝ=��ʍl������Q#^���}O�"��Fw����ʽi!)退�mmN�PJ��R��Y�ڤg����)�=�t�9��a�?��q5�m���p�'�o��b0��:�%I�J�H��K�Y����������j���t�Q�hw�S���Z�S�O�������C�r[�C����S�u�c�䯶�.=q��Ŏ^�YC�ֱ�_�:[ó�Nr��x�q�wG�5"�W�#�uB�@;6�q���D%���yܣ����WP���V7��&����2\�ać�I�Jtc�H�!s��GO&R�ga��^��I0-N��v���"��Z��`P@��r+9"�j�˪>G�5�%'ccS�k��_�߳�;3솿|%#P+���Ҽ�c8�"^��`�����7�\\v��'M��x&Hڏ�`�떃��g�KD��Ɋ�9�L���V���E�
������/����9���ד�QR�	�A�^"G'���-u���55@��m�Щ@H#����Z|�Z"F��]�i�{L@��n�~�:�7��U:�L��u1���7�v��*Ke��ܾ�3��d�I��7B��ʳ΋�/��]���ibލ�]=|�ZSDN���$���Hv��:����+3f2-�*�r ��&���g��8	�"y;tLn��/!�k�jjy���(5Ő��%�9EEAM_���9��xk^p�=����!�����<���wk}�K��L���p�L7n7�v���<7H{ t��}�@c2��7����U'� �<�F}`���,���ra�$QI���H�Oii.~s��d����A�m�[4I1��!����lg���v.��
˝+����d���`}4���|��i�����
����Z�;%�ؚ{���";%�,�p�c7ji��飦��E��?�ܽ��S�0�>�Pn �:͞�i�L�ó鬩(�7��� ڥi�g��3B;d�g%aFj��GzS�[`ST�X"����,�����L�Ga�T��;��I��3ҝ� W/�=�"��@�ʰ���,�f��˷ �x�G�,ard*����8�L��=�}E6~\�$��uy�	x�A9v�'R���F����%�� MZoul��=mW��*N`��{�L.^�Uj�[��Gnk�!�$	fil'���AH����y��	��2G�>��e��en���:F�#0�B����r�R,�	�bf��v�7��(;�D�ou�tВ��!/��(�J5r@Mv���G�7}A����7���3��h`�ޙ���`��Z�y��/׏={w���>$��]��/Q�8�Oz܏����_�q���mF~�~�}|c�9=�.;A��F�ޢ��fZqi�W��[I�ܯFdLF��ҵ�������K�<�đo��G@'L+͟|)%�������9��/����T�n0g>E��GX�Z�Z�b�Omb2c+3J�F�*����B��H��4}9���5�I��x�	�3�a��
�n����b=?��3�z����� ��t�0˓R�e��cj���s�x��|D�����0×� �`��*7$��m5~C���m%�4&�].D���6�� ����z����T�*rܖ�Q��W��jՆv%=Cp�nP��~��[���h���5��:֙����="��T����0iާݣ�~�9�N[���<���}u��[��7��Ѧ�H��+��"��=���_?�l����)g��R��r�S�/�#��d���pK��ɺ�
��"���H���+�(�6%=&9pw�
_��pgc�kli�d���&2����}"�!#�S�Lb��몜	��]��$��G~*�����\��E��quڈIχF�:(wƝ���	�\�=�u*"����?�<f�	1
�]h��Z�ۮ�j4�^�J2�L#��4�ʳ�5��CJoYS�P�xqj��ʎ�_`�L�T\H6�nI�1�υ��^�~�Fz�-"Ngޅ��l����ӖK{�h�`���o`���‭��9W�[��?����Q�]�;J{
�r��󻯮��y�g �^Y_`%}�9e���y����P�qKR_!]E����,?{�5��� _GR��;l7�Nv�e~�zHa��|��G��j���B	�~PCc�GPxO��Qo��hȃKH�z	�s�B���E((ڤ�݈��������t9�k�� ����U�$F��橜��:�g.&�b�g����;�Q`=י5XZ��G2�2���ڋځ��~ۆ�|��c��",Ť�,�'��Λ��[0�t�$��*�|��-�&'���<zw�mc�֌J��Τ!���,6S��%�ۥ�b�qT�JW�.���\�!�� ��۠ni���ƕ9�	#�ބSs��5�Ŀ��k����ɫx���R?�TZs�r:��&��]S������D-��}MOdR�)-J�gE�NŢ�C�p��`���4���K��-���+g�7kF7��K㵾J��uū<ޓ2�Ӹ
Г� �:�[zH�i)k6�v�?�#q�G�M�Q�:�����r$~�B���%������t҇�4���t"
q�U�)�E�3Ũ�uΫ��]tOz�r�V�68�7+d'�I~����Ʒ,)�ST��ou��Fñ��xK}�z�Ov���ф����D��!�w~޻�w�6���h�T��l+xN���S�C���
����B�fW�
|�[u��&���k:Q�1�ڎ�L����Eu"����%��\�8������/y���<C�8���(h��C�n�n�n"z���	�mSZ������[�p,�W�$�򹷰���*�J�Oj�A�c��<u?�{[���s4�
i��ucF�@�j.�������XgC�^r�����u��B]�0�&V},ɿ�x�f捐� a}f9��2̡3*te�=�r��	2���0�|���7�W�P�=үZA�� *�sI�KRZObu�G���Y�VBbI��i!���Î#
^�!=���
-b�57D�W�|B�D2�p��ج�?���*"��G��B�ّ���kW���,���{����F�z����l���i��`�
 �r�m��v*J�L�ᶱ֢.��u��,_�/��ۡj�n���)�U���q�ߔ���6-���	�ѿ���ak�9�a�C�(��T�����v[Qm���Ga�C��΃-X�%`n}������f�@�k�ŝ���YVG�	r������ ��O�e�l��������d�%1j�%�<����<�����Ү]��lgJEDW#����V/-|������`ɹ����e��oƩ�Z����o^[�?�����{{�e���{}�����sϗ�rv�K�PF�>.1K��x*T�����^J��L�}���g���)��<�F%X=���E�6��Bbd�e�D��!�.����{������n7iV i!�N��@�
���MMH��~E} ��/2B�![MJ�E��`׳��9ɫy/�R
ҿUO?���{��d�SiJ���KPA��y�b:Y����o�4 �/$g���~u*�aE^{�t��ԏy6x������4lԥ�h{s�r@�J�67�E{iX�t䨑4֟f�����$�e�ߗș������0�VD8�=X� ���:@o��&.mk�Me�{i����w�6w!PrZ��9����Đ���
Ng~?q�l]�����.��!�3@JC���{X�9�Z���U���&�%��vlQ�KP�\�Y�_ c�)�6�%��A_�(P�k꾬;��D�Oz�nI��[�k�e�@ ��mm(�����[��z2

o�tӯ,��B�t��Mv�Y��6|gq�{�:����ו�*�&�I��[&����Ɗ����)�Uk0��%�h?����Q��'P��z"�8ڸO��'�� H���^��X��V���l��d���ĐX��"g����?v �$R�}�NǾ�Q�f@;n�te���,\��xB��2�@�XuEւ�Z�Q�)�fһ�ʡ�dD={��nA��I���Z~���O���V4}��_~ئ�!q%d�{�Iv$��[�O��.��áwV�HX [S���ˀ��'C�ǞI�(e����W�m�I(�[���$��4�z�x��������$!-�N�ző}��,�b����f�,7�U��y��}���Ƥ�<���h>�� �����=Uk��څ{~;��>Z�}<F$_1 `�%̔������L��/b� �E(?�ĳ��MP+h�A��(rQ�>O�N���3~����L��q�f,!/y�L��I�8��J�L^$?sK�6��)�|'܈���-7��|�l�,=)��i���p�?�$� ��`��a�xo(!�[�>��r�^��z�u.QG�?47��r��CD�R�"�u�$�܋�ɺUA�I�"c_γ��6b7*�L������X�:��y@�J �ZԲJ�Mm��y"��]KS�'<U� oz����5$�5h��З�E)a�ND���e�G��CwJ�i*uA5��v�6$��aa ���iF�-(;�pȟ!�d+�j%�5m�)!�c6	��,�X,nP����TҎ�G/���5K���K�3Q�1�}pT_�(��r�S���f���U�&^'cY+%m�
H*��%��{\��C�T�Y���G������	��=d9�2�9@lq���%��mw�����dv���b�
j���;1��c`��g��f��L�t*u-��PQ_D�Kw%�C����J!�c:z��Rv�wb@��._(��M�߷�5��)pؓW�|L����#'�A��]�:�D�6}W\��|�"1�K�m�o$5h�â�d�D!���j	��U��!z<��>�wO�E��b�t6 oBC�g��s��?b��Ii�Q�3�~��K�;j�k��%0&�(��܋����ƅ��{�������Q;��-i_�&�v���	�C�4t��8�,����H�R�1�/�����B�5��5^�"6!Y
����͵���%�,A��/��L���i�d��ۭо4�����Q�w1�)�3�&��~{�'˨��LH�ߒY}�=С.[K����K� HP3t4�f�N�/�<��O�ۈ�,�FEGz��g?.H��Fv�=�V�؟�[�f;�%zkں�F�r���*�Z�x����-�OꀹQ�g�F0���W�������C_z���r���C���@q��Nߍ�*Lw�H2�T�ژa���\��,I���wGR�DF����2�0T�]�,V�v2d�_9���N2��pIV���oN�=��t�b7D��bE�t蓘� �V��!�8�%
�?͔+��"n�v'��G偭�=cb�޿Ί��=���x��l�"���Uw4��ݼ�<2�����5{Mm���L��)�&�a�#W�7}5�fblD��������;b�%g�\��'��uc�Z9~�hv���ɮ�}����xUo�V�]dF�����Q)�{b��̋0��#�*0�<�wD�������I'����T�3y3��.X��/�B1���{�=�<�b�����A'��������@-4��o��Ӓ*&�����-�>q��`��퍂�I�(Ϝ�=�L�q�}�Z�.vy�ӗT3]���>�K�|^�BSQ"#	$k�]�G}5���XN�W�MG��� �?"J����y�R��k>b�����܋�P��R�!{��γ9��n�wى�pky@�K�{����h���h��E���2!��l����k�⸧�h�?�Wq����^�D�j�/X�ͅ#ST� ��Zgl0�L������B0�z����%���c��Pk$_�B� �~����,��^OŖθ�	�۔�N��j�cY�d7�|��^֝�Z���������8P��/�$'c6ɕm0�P�0�k�|'��7���Y�>�%�=&�K8A�v�6O�T_��[b	���+a����D^�
G.���	��������
+�L���xɷ��UU路�v��M���v?�7��������S����m�To&􇱯*4�����AS��	#% H��ve.7P{�yD0AMʝ8�f���V�bMޔ��L���$��gZb"7��� �u�;�0��|�,"k��ΐ9��� )�k�Ph�y��'B�jゼ�[���_���n+�>y>�y/�}�:{#�2��Vݶ�+�|w��2���Â������	�F����{{O	�2�Z��}(���%��%d��������в����;��kP@�S����ÿ"�*��΋�x��=� ;S
M�P�4��S3�����61��P��ي�'\E�k�;E�[&��k*`50�����9�T��d݌Qi��3�.��ķ���զ�PT�i�O&� �P��E�����,G%eb��9��/��%��z�����Ñ}���lgy���X���V�g�^T7�_�M�kr5� ��.t�BiN������i�ni�L<j���@��}�=�8����2A��䛯$�O5���T�Qg+j�x@<I2��-(a�g��FK�ʚZ�瘥寧�.i��z�����:�E��3f��>��1Wg����=Oa�y���'8K�Zj?�CeS�F�cgƮ΃��#A����ZL_1��9���V��m�}���e� J���������M�����m-�wԒ_��m� h�wv�·�m�`VT��/"�T���G�"xʿ0|a�Wt1��<���m�g����*����D�u8��ܒa<��*șM7�c�Kc�����H���5*�^:������\�'ך��|�r�����o�ڨ-tHs�Y�E�|1�{,l��^����vF�^��က���vM!~�̪�-	��)0�#�� u�p?N�f@R:�ӳ��aE��c�.�2@�$�����S�!�2��n�=�_�;$���"bU�f9;�ϯ��JcÑ}�I��(��8���<��.BD��@�p.��M�FZ�#����n��Р.�)��قշ��A�I��3;�x�*����oƯ)����PRڿ$̅M\���-\T��ȝ'���š����0��$,��EC�6��M�+3�\����{�ȍi6�������{2-�����#�����ښ.l!��S�Be�}�ʿ7ڒ�)��`�杈^yK�z��i�iF����ͫ �?{�V>�G�c4b�(�v���`Y���Dg��MpF�lA�!�/�+1z;&��3I~��w$�U�.�)�N�O� @	e8��� �@4Յċ��V|$|������b��µAe&$Y`�_��`�6B]��w6��U�ܧ���Zj��dLr|P�xl�")�jbŗ�-㩰Y��4��A�Q�"fD;!�g����9W �/���[�":��Z���+�&�����].��0��0�'9��;%@���p�*t�2鿺@��}��{��+ot��8��<w�a6����Bh1���{ �S9x�4�*
TR��Fmж��6����L&�/�1�Qg�ea�M�������.p��#t�z����Z�n�;�^�{DX����x;��)�i&�D��z�sՃZ�YJ=b�&N m�%�
�d����]������3��:�F�-;�d�sk���l�꽮� �{���c��'�������r�7��k�	�KJ53C��wNO`s!%k�B��������r���{�k
�?��]:�d�5wԔ���ŷo�:�fZ� " VV��Q�F|���қv֗$�Q]��P���n�R���9"������Q��q=���\]�a��[win�����'LMq`��)*g��3�0��n������.Ug��Z�6\4����Q`�q��=/x�˸�Q��(��5�m�FZU��۾$1 7��A )���s�(�*}�ؐ��=u!�)�!��[o�`:Q��l����,�N�h#pN��YJ��^z�؋v��"�-S.���±'�����L�Lp�M�6t�hN�tU�}���C�Ч[�{����� �+ ;QHwR Ic-�"D=��`���1V8�Q3�M2@�*U<XC��i���CcϏKۤ=B1u�I�J��0(�7R+����2��B��5E�i��Q��Ԇ��#�ܝ��;��`��
%|��ԙ�����3ZV�q8���^$")B�,K���.�e/Tڴf:�T��&|�LV0eR��F��*�~d�	~���*!�t��vv˦�pNY��4��X�:	�j��CE~��w����Q���+��b#PM�p�Xj���}�*��^
�R��K-�d^�����s��]��=\)`1����h�yb�@�������/�`�f\�N��y�H�[<�9?Q^��)�逛���;�*��wY�\}��}����ñ$���t��XW���[ў��$��;Hg%���;"*���)��Q�T��?/ZJc���$��c�M8� i�aՋ�Ey�p&ʗ�F�*���6 �QPC�י@^�R��zt)���a1���<y 6�+�o�xR����%�v����D[�t~
9eb���{</ zH]�{eu�)���*���L>ԮX2�0�l|n��]�[:����6����"0��xRc�C݉ϭ�Ք0LG:���}�9�Σ͝���P@<�����Z��2}�c&-���B~�i\�Y'ִ/���"u�3eK�2Y9��dTv�,�J�0��o� ʲ��B�}�I~p/2H�/�MS��v�gm������{�cg�LK]����M2"�D*rF$M)�6���:�Q}�c�e�ps��@�-9�Z1��A�*g�d��2i5 7�d��*��.�7eYzi�7�5��q���y�<ݼ1x��/�~
�>���@q�U1_bW;��' ���Ĝ�}��s��/0�6.��g�k��m���:��t������I��:���$�J�[.S戛g>J ��b��"�P�	r8�NUj�(x#��
R�]�EWH[�G,��f��M
-���f\�����dá%*I���V� ���t�4��x�wJ��}�ʛ*��{Q�Y�JY[(������7�N�h�a�����
�^�m��]x�VLnu�SZZ6�}�>�OAڰ��S#��.�-��k�#�t�Rk�c�N�U�=���·A_�븟ڠ�N��2�eo�'�Wu���x9j���\-��-uji���D�����cWE5q~�O�r`%Y3Q"ōlT.�1Y����h��zNLIX� ��ŬM3�5`�N�}�mG��[~n~�\���t� ����l�ӥ��9N?`����}���άE\��f��^�N���.t}65��|�TA=�Ȝ�	�����΍�+G[���{���-�Z oت5����j����Xv].�!vW��R�>f�1�;;5��w�L�t�u-�B��M���m�r��u'��zP��C1��D:�Ǩ?��v*v�u�C���N�Ĵ:JZaL^yѯTc�y]'��:�|��xRd��$/�:���g=��2ER�+hU+��A�p#mK8�0��<��<]1�{���'��?�M�='P	Q��⛝%\���F��jX��n+��in��2̇i�Iw�>a�\�%�^�����N*?-v�rS�\��f���P&�F�N]��Bp�M,��a;p�k����=�q@Ļ�@���ˡ��S$���������0%I�E�!��
g?������#�VF��.u���2��}��V����������S�1h�/�4�~,����wy�[�gX�sR��� m4��/�Gn�.gj�I�G�Л��0vű�O�o�Z^TvϥS#1:�~&��H�O��5H�ť�tRHʾ�p,�'K�<u[K*I�=]ӷ|=P!�m=#���t�nUa@�(9�>�b���.O��#� H����0ż�Z����3K�����;zpw��]�r��.�+g�{�L�³t,4Ra�z&]8P	uAօ��m�`I[�`IU�葁P'�xg�!k��(k���uD���S֟��O�q�	AΜ��0O��ݶFq�04[Q�vټ�J�#�����os�A\�x�����<��J���]Ncl�g�i �����Q���E[L��"C�HQ��GG1�3��} TtlN������M�7��l��[i�AeYܽM� �{�e�5&ʈ%�<B���◱����l�HDӃ]x��d����K��uO'��oT�=�*����$����*|�U��t�s���Zڧ��x2��}Q����]�g��z��>=�������,hq�?P���0�؂�L�2�<s��{!�|ZC�����~W(.^%l,.3��N	�S�0�G 
Z9���_y�b�f#>�4����������
� ���	.�gBET��Z��9�d0�!j͛{t4�̔�a���H,�[�||���jt� �n��y�����R>S挅�i_36FWd�K	�$�"���5_���05������b�KA#�����Pv@<�uH�����0s<��So q-o�)ۜ�J�����Û��<q
��K���S�9��v��Y
��Q�*	j|�Cu�j�X(��n:ڞڬr��s��A�!�|ƌ�(~�o�^>}:<�+=����r��@B� `��?�ܖĶ�:wJ�r��&�7Lc���Q5|K܈�D�{�E{�Y'MFe�z��A�(�e�1Ҁ�X�n��� ���w��h��S���4x�ľC�z=����o��<|@ܣE�)�
-fwR8}���N[ ��6b�f���tṀ
�Ld�=!��t������a/�6���E %w`��7CICm�}��r��~��'8�v���&�]���*��e��d'�l!J�4�"�z
�I\�=��ؚz��y����)F�-�;�)�`!���M$�2��S`Z��==E���@��[��/xH���N�\vK(o:}���RK-�/����AC��Cl�a�j	k���R(�U�3f^��)x��ZF� '��¦I��P�cS�����^�*��2+���-W��x.��*�X�^A��@���/L�	���=捹�r�����n�3�}����buu����?fe�Q�7��x����z�߅�p]���V4s�|��qߖ7OӼpF�bA3�%m�oaި7�47Di���{�7��.r8�ꎞn5I~:H�I3�~NRȈ���R��ĭ���1N�;��}�;mU�xT��-���a��A��T�=�ִ�O�?e^'�u�8
e2��zUdh7T�0KAL+� �~��5 d��gJ���lP�t�ѿ]dn����~��XM�x�3&�k����4��}�= !@^��/�Y�\ r��uY�#ry�Qt��1�E)7�6�p�71�����.,���l���^�	&���6��N�~���q�q�૴7����%b��.Y_[�~|�7�l�F��ܟ�og�JW�o������hqI�5'�:o,Su�)%��v|��f�{<^{� x�/� d�R��n�-$s�-ģ$-��4⌷���I�L�o�{��3�a�YX5���,��;��[Ąl�;��!5���9 �;��j���� #�d��/���'�X��I�D �۰�����
f��g��8����qn�R�z��]�XQ�-�ͫm}ٍ&YJf�YsR�oI�C�B}�UZr�iN^xCķB5�!�l��7GȮ��~����}��<u�����zb3�)����2�b�GK�j���������g����^E�n�� `"��+s� ��T��[2�lyU�� (��L����w�N:��=�"�2�����t�sô���]�#`K>��w]X�c�>�@�����(�����q�j�KF9$�,��5�F,fp%���f��vֆ?��W�(t ����O�\���fUe
~"�$��0)�Z�F��,�s��������Ҙ*f7���X4�=)�H����UH���w���PQ��H�Ɯ����(^5�RJd�^��#d����` XZiv����^�3�;�@�z�ȗ�x�ں�V�]ɏ�t��zh~����]GS>Ox�5d !��"��^��Q�~l��~�,��V�0<�
׳Kr�xuW��䫻��U��u.�� W]EՊ"S�)��}3h�ag��S�t�c��A�*~x������'��0y�i��c��+��U�fj�X��UT>���-!�c�z��=�~�a�*uy�<&h�&�,P�H�V)�\�w��L��%`R������\iHO�����Y{�c�bH�J�&�(qj��w&\.�+�p��������V���b0�}0�|���*W���{rit��%_*/�]��Ór7�H�����޵~�e�����H��˅��ҏ���b��얄����{��4B �{�N:�����:z?PS+GG���L���|吖o����'�K�㻅�I�[�t��i �o�S;�X�[���!ʱ���46*c�4=����ꍵ3QD_��?Oð���El�sD\A�1Aq$�y��2�9ʞ��R���Y�����q	�u���;���
FM4�l��mr�y\��!T
ݝgV.�w	??��K�;�p.�^C|x�\(�3�~[�B6	�թ��c�߯�h�b{��4N#^`"����Is~w .���~ %ya�>���m�N�H��,��|��汯ٴ�,D�N��:�_��mRUO���J�pg�G
��W�HC�)�qiة�h3��l�H��i��VHOҠ�Q�"��)oy3dDP\>�̾������hd2��51���=����A�;]�pu�{�~��Av�/(Np~�eV�7�E��
�q��'����(¶*~9��o#��^����[�� 0-��L*�y�ݸFV�~�'f!;�ԵI3o������������� FQNb-Uv"���}�/%w6c��hm:T��r��.��$!�7�{ċ����oE?��Vé���Cfq���J�&��j:b�H��G�Կ��F��ZBM�V�0׵0x?Y��9������_���t��H� Ú�G
�2�~y������|'�-l���T�����U�D�mJ��)�FAYL]�������{j�QpH��Zԙt4�/�DH� �Bp�n��jh��VJ��?��a��EOᗰ5|/��?����\R�1,��@�mHIҪ�M�vt�i���k@�ч��8����76�Pa�4h�B���ڜ�?j@�=��õzl$(�څً�i��������s4��^�h*�נU̷}�i� �[���j����5�c�XR�a�}S���$�{�Yu^�p7�;��ҹx-:�KG�|��G���s՟WO�	6��[�i�����0ߗ��2DL1�.�k��v�3��;\P�0e~�%�B��F��>�
���V�=܈\`~��ίE���Iy������D�q��D�I p����J����m�������~8�P�e�a�"��&���.%�b)L\�#(K���`��:�[ث1�h���ɜ&���o~wǄ}��c��}��MW6�����&(G���A�U�������)m��.f��%�{�TVF"���?���w�,عN�R��GC#6�W*��~|��x'�B��p6�|ʱ6�=�6ē@ ���Wwh����}��=P��Gm�5fms�{�OK?�4����u�t���_��ZYO-�l%D��*H�"0.d�VL���|'P,�	��'o�ې���W�qO�;ù���
�+~X���1f���+�Q��w�?���&���d�	�?
����������>cbBw�C��kP�N���N�hW�"X���qe�lp������u�@��ʌupe?��s�j|s����%�A����7���a�c�'�8�K��	�_zV�������W�L�G�=�]x�p��8:xl�F"N��!�xY��z�9�<�ҍ�>�N���E�� gO4��5P$�O(&Cr��=���M`�	|�V�.�bj��>���a����d��������0�_�z�Y��iD�*�I��ƥ�
�aa*�3�*�J�,�ړ��7���ln;8�!�c��E͜�]+o!�׹=�"�_�A;�%��JL�Kb�lHUW-�:�y�OU�3[<(8�Kr�� 06��Y�����8�\61��J���N&��e�T���{�������V��p�~��`��s1*���q�T=Z�h��¶~���a�<����H���6�=\��w�����9�/���@�U��엺u&��v�zx�&�T�̾t��c�����}�"���w|��|>���#���\���ۊdR��x�'����+j"�Kݵ��2;(4�hc� �s��0��yӋ�]�g��L��Z�?��!�]p���ё���nԼ��{uw���1 �$�s�oI<f*���(pL�9�yIJ6}�n���"#Jf�D5����R�($����������8���!�:Q�0]�av^	�_�?>?�G����ȷ3�k��*M�b�p�	�~�"������)y����7�5SR��I��Ey���&����?�{u �O}�~2�0�<H$��O�Y����L��6��^"|i+�S�B^Ҵ��n�I�h�!δ.O)�-"Ng�n'�c���Bth������1�T�� �R��T���?�f+�@��C^��.�5�8}D=�o�1�h�Aژ�ӟD3ƙ ˿���A!���C���%��TeT�\�� ���։L�F54)���nq�ܑ�$֡�_ i�®��v�s���k��쏈&���X/�S�N��᫨oR��7��Ю�Z��)����|�6C��ޞ�в;��u�8��t��KH7*%T[:�n%ھR{�A	�t�H���.�XjR�O$9=��V.�ſQ�s��`iY:�>`xT�j�ě]z���&��e�b�Ae<��p��4<�OnT��O�Q1;���܁B���ji����e�b@S�/r��P�>��M��0����lH^�Osz)�F�m��L<��']B�����`���[�uuT�=T=��#�"F
�z{��1W��x����ԼG��+�w�?q(
2T��4 ��wp�������Җ¨��޵lٞ8�hH��
��6`���XV䤴�dNB�4�h_�a`hn��~y�\��+Ǘd����(�u�l ��*��
�f�S�Y|�����i�4ݡ�`:`ev
֠�6�i�Uby����[)@1���S�ᨁp"�����OX�~��|���Zn�yCj-[��#�\H�2e϶f���y����;��ȃ��EH �ߙ(����<Vؠ���v)�0��>ʑ���|�E����h3�;gk�o�i����%��l���x	�Z"�\�����E��B<�b W~~��HM"�U+�ժ��%���^�D�|{89�ʥ�.}�S�7���V�	F���|E���́b�V�yf�,g�gv���ȏt����3<�ˁ�}�>i���?	>8���t�́�ty����4�����*�@��<�<����3� PV��z)��Kn8Q�V�Q+�hu`
��%Jw��>z:��[�I��k�
A�(��2�A������:"&��p&���
��%���.�]��غ�Nm�n$9�M���j�Q ͣ$u��n$����R�w����M�g�2�&������1e�`F�a.����p�s�фhrk�@m �t�B��,9�@��"!�3|�~��e 3���R.����7����?�ѥS���G�7+��4������I�w�U ����J�\���S��!���`_�\>}%:�\J�}J���K��W�N-G��=�~��� #������(�*[�,�oL��tԝ4D��U�vy���L�Ʊ78�9, ��O�쵮�^��Ω'���дH7Ĉ�o�9��'��1�ݹ���D��vy������V�j���hv����+�_�%�Y7�����i��\��-$�x�)�{R����P@����P���5�xOaj ���-��bu<B��t�	�[C��K�(FF�2�*�+C�U�4U<��8�ح��2��$͏�	�/�tǁ����Ҳ�K�"��I��DT��?��\���|*�A���42j��C�uC-�[|c��$'P��?e�n�jفEU;�Dg���K��-qa�?�ڑ��W9�����t`��'nn��'�01�ӿ�Ae{Г���1��� ;�i�墉L��>��~��c�<ȗ������;��.��3,�B\���^�x6P�.��D���P��|�w<�Ζ>P�?q��:O��7T\k"�3��qkzcp��Pɧ6���A�F��"����T���ը�$w �;���ۜ�C�%��^���(���<'D�]�%���`�ڜ���'|�=q
�4��S}/�g��@��u�k,[Gr�Yu��͟�H��d�c�%K�7��DӤ�\[?_���M��_��Fv����W�BM�!�a�*���Z����6�"=�?��R�-�>�h���=�B�/���>��Y)�,:�e0'�]=�i�ST��;cb_���U�"{���e�<Bq���v8���5�1�8m<�ہY�M�;�N\*�YƖ哈��Qq�F�~�.gE�~�(�U���n
p���2�)��0��Ԣ��jG��Ƞ ���b�k %_�"rgW
f'��
t}�`��CGA���'68�g���l7�f0Ǿ�py��7CPqH�B��""���M'�6�5�\�'
t���C��p����]�p�N�ũ�ل���k�_�u|��	�L�?�˓���I�6�p�hk�l.ɴBr<50��к[����K������!e^ǖt^R$�@b?x5E8����h�o�EZ�H��z��=]�x�N�W@@@��k]��l�+���Q��Λ���7�+D���1^뢉8|*�隲�]l�^D�z�5�W'*�����|г�������'���(	M���z��.�E蚘���x[�6�\��=�S�Q|:F��9��4�p����C��y
���R���P������BY{�b�e B*��u�j{�{�M�=�Q�p�C�#��9�KB�3=��m;�n}�.�&+4��7��d]�ɮ�;�E��R�dޤ��1��񲿃{���l9as"�������W 3x\�<�X���#� ��p��n��ϑ�K�9�b�Ȝ1�r\d+&�;O)C�C(�4Zʰ)��~Qݡ�#��OC�������W;k���P���xaM�g�?�?�@ ֔P�P�����Bv)X����w���ojnK��i ���\һ5�
Q��T-�<U��9-�1d���'�.�H�2@�����{�Da<%p�ބb��o����>%����x^G;�^7@�]�[��DERì�p���P�����f�jh�x����+�E��H�xc��C#��٩�65�I!:�Z���'Rkw����費�6���@���������NĖq��U�ca��C� ^)���]�;TˮO�9,pI�PQn	 g�n����8��9�a#��j����á2�c�8�ZOPmޞ���q3��ӳ�����)(5՞T��>��x�3�� 	�m�:��c�8���r�hWf9�T���B�ؕ��ؾ��l�m����� {V
z�@U�My�~���r%3 ��ŜOb�'&�`�F|�(B�
/a��w��NOذR��^~R��A6vÊ�*���Q��N�Xa�a��d����P���*�[����h�T�'�i* ���y�@o	��e�p~�i�d��d�x�^J��M�#���놪����2�p�ݤ܉�G�q��č�b��	�`��i��j8��og���gG����Q�^��y���_*֦��r��J3@�.�=�HO�0Y��V�k$T����*��&4��Ӹ֊�N�W}@�3N��U;<�F�S�_u��JN�,^�(�A��!?�Z����i'@K�q����W�����]���$DWqJ��G�5p�7�+\��4�˜��-��9�h�)y�S�Q��l{�\HH��*�e���MK��Q\�_{��D�/!}���8�q1��R���W�����¿!@����F�&X��������RrA �R�6��ۡK2���{�5�Hh�H��,\��le�>zc��W5��8��� 4�dk���H5rɀ�;1��<U	3N�TϚd�t��Wf���b��H��kz��rӳ�Ɔ1f� =?������ [������DKg��-E��I��,�nn�^)�`��b�}���/fDS�T����ǚ��Z���=�Wz��B����"���p�L����J��!iS\{z?v�O�NΐI��)����� "�Ҵ}�Zw�-��_�k���ـ�r�~lWe�tQP��y1�0&H-$��'���"E�U�"�F��{�<�wB`�Y��q��I U�K���k�uū�Ĕxv*��dāȎ¨9i�adĿ�@�Ӟ��F���
��D�pS��C���pN������Q�nӀ�+r���|I��� �U۲m��#��i�<D��9jXN��^�n���G�Pw	�g��Bٍ珷���9�1Ǒ��W��*d>��B�B��T+�'ʻ������]cɈ��X�PI����ͺ���+��w�����Sh=*����H���w�:������Ẉ��$�c����_��]�'���֍K�����}	�*(��	�	�.Mb��f������'5�f���Z�[�NG�'��,�wM�դ3��UB~^�7�"���'.�0�bZį�I�g^5 ��N�����Js��CR����Q֓]z雷�?�N��J~��e���ڦ��F�^\1�ŀi��N�4�x�~�j5KJ�̋Cr֏{{BF&��$_D]D ���H��0��s��?P����듒�����Uu݇$�~G�����Ƶ2!�`�!<�� ����( oR��,{~P��OG+dxs�H�Ya��z���/��*���Z��e2Îm�M�.�~�YǄn$�ϩáxWn���L�u �6����nJ��s��+ �,U��@�7�t0TnP�?�a	�t�����P�r�s��U�L2~Dq�lQƾ4#j���~ף�tس�-�ǮeY|�<���˴r�-��:��ه^��&�8lP<��a񗥰b�h��o�*>�s��(�YI�.��l^�Ѵp��5V�z�aTnuz��s�f0*��[�6��/��RR�?uc5��)ݻ^�Tm7!����!�Z���@����9%z<.��^!������V�n\�*����D�k���~)l�ee�]!�g(X�+&�KF�E�*��9��( �����2�È1�]C���i]���8��	Z�޶��z�6�����d�1ɸu��3�����+z(@�
(�hs�>B$4w[ts��Wz^��D��OK�e�Y���f��^C� 7�왆�e��Z�{Y=���=�B�����k(�\��|�9��V���neH��Z��Fg9f���an��7B9`0��������l��F�����)�nIp/�סx2�@J*o��}q�݉�M9�\đcc��;�M��ȥ=�����pp�)���-�@��8���~��0����د�k�p_n��Fs/`�i�e� ZE��|m��a��Ϩ���޲A+F$R�w�׊ҫ)�o�#.�h�7D穜Ȫзv!�]&�o (杉���ޱ��X���;&�	��+�����0��w.h�4[��%'�vk���F,���z.��d��Qq���C�����j��ٮ.h��oX�� <|�<4�t���b�oJ���I��JgDˠ��Bz�́���ݣ6|�8c�9��hNP,{��i��U�\3fS���xs�$�Z+�;�Nf��{uKѨ�N���)�L���9vO%^��a��o�� [���Wݤ5x�����7��i�)j����}SKXi��e"5ܬ�8K@�7T�	ѹ�S�w�+$ei�ÙVK��h/��"VO�A��r����*��ߦ����&��������E������:��xQ�g0��7"�>���2�_n\����@g��[�Wm�{�c�Qju�i�qݞb���b�ʉ�g�Rғ[8��I��پ��N�9n'^�UB�Ċ�V} ��(�<�;�*ov��%;�xX.B����4�(Q.}�7�c��~�Ղ!�o�G��ʭw�x��ܒ�C�c%��#I<u��=��K�����ƦT��t=���
{�sVhe^�ֹ�jY_�m��.��4�R�9uAk+v�T!Ȉ�F��%��L�}��O�
Q�:{`YVCW��]����K�����lڵwv�6v��d�\��3���ޛ�
l����U&	���~�o���F-�^��[��sKJ��Y6,�9����;v ~з��Y�8���6e�[/������-5'���'ƀ��]C��6�N��r��}�ؖb9�]\:Ev��`�tz;Z�tS�%Q�tb͞lN��*\d���
��n3�hT��׼��8��ʩ���Q��0h�][Zp�q�b��uLs����r��/���	��'�E�|�?�-q��Cz[.�)��W@-�B�: ���$����4ĝ,�Bwx�u�GD�*Nݱn��x��p_q��=�WL�ڷ�����\�����ʁZљy�C;��$�]�&��F<#ݼ���-���	�u@·s A��Y5�፪%@�0�iշ��>��ɥnD��WAKw2	vV	�w�d��z�����@�"���N�����ѥ>�����_V�|t~
Fi-aF�:{�� a̻�MH�z{��vq�P��ƆQ&y2��/��1rc�)͗_�9>��4c�����W@��բC��A)J� �@�^9���P�틊�����B^��j�~ö+����	��7o0
*�����`��Ѷ��r7~r�-ݿ�{vo{:��5&�To+M���c)%yMN�����/��Io���b; ��`�Q0 cw,�Q�9�d(3A�gx�p�/A��v����'�?86XH�� y�kR4tĭ�`��O\mHs`^�S�������N>������z��F�ò���6��t��G�H����L���d��)�~�F�7A:�5���Z~|���mfa�~e/�ۨ��%�@,폇X7�����tW��c�q��PO۳L��iV(�{�e��(��-���-���Ձ���`�hªϋ�Z�zEub h�$�O{�}	J�͚�+G72�-`��~�����<q+�m���4�2۴�nr$�V�Ư�;K�M��e���З�0Q
WhLmI(BВ�P�v]�_�%['{���)2�坴ړ!��c�"��������ʭ\I�[�0�/y�Iq3�[no�6�#P�4_��X?Ѝ�	�2{l��`hc�%0EiP��ۄ�c�.���75	�O�l�[��uJ�!f o�Z<2.�9��h|
՞�j�=I~� �u65�(�7nU�����E��(�?�&g!#@��G��3�\�μN. s.R��ʦ�ꫵo�5fc{a�Y�!��[ܧ��Ӎ<�\&����ȓa7$Yz(5CazD���p�t4��e�S��j����H�4A�vZ��^V��T�.J�`��ֹEI޶,@��mj��Ș��X7#��O,�8:�&
���R�d�#��ƻ �x}��ɫub|��ã�a�[#�&	�E�{?��?e�㇭�f0��� ��y#�`I��j��?�S�e?����:�n<)��H�̂�+ݴb�Fu�~����=��ڒt@��Zhoٽ�����ڷ�gK������N<������W���6�'�F�����tT���J�p.� vW�V��4+R�6�2���ayȔ=�p^Z�P�e�!v��\{��a/)���7����4'@��]�&T����>��kU����D�[�b$��
���#Z����s4<�=|�G�j��hǖ�v���n xo����M��;�T6��4�R��M��/例�)�G$)�pԪ�Y��Z6M���s����A��m;�X�d_�N
# ��S�iqT9�����ޛ89���K�$�*/K�Fĩ��N���sqc�M4�Z5��:�k�L�u�g�̢��!h/m�l�.�C7��SK_G��b:��|Ő�xk���ihrS��ͷJu���ʊ�"�#��C�`�#�g�����5�W?�:ʣ�=-��E��UXޮ|�Ď\"C���mL ()��L�6�BR4@ٳ�U�TXW�M�BF��O�(��{Z��t��d���)����2�x���S�S�;BK�28S�n�I���<8��K6^ 5��< �9��_D;g��[��i.�=��m�9�3g_��B�pz��qG����}���L�0n��㚬m��Zۧ"
3Ѷ�����F��Wq�U=�
�=1���{d����4��l<!v�Fq�׌�^�j�V�w`^�rH�͠�Y�A�^��E[_����~B�g�D���m����@�>�I�0L�)|E��K�9����;|��0�WJWQq��T�7�)2���r�+Tv�!Ε՚_8�;�aB<����S�a��_����rş�r_���b������pH���C���+��.d]�b�)��L%k����rM��d��5�h�Ö�'`<���z�
%��l7 Od$�gA����Zg'��M��C�KſІ�t��c�n-8tZz�ԧ�$ƺ����ی�g	T�d�G�-�T�at��F�2�Ռ��k�Z?C�q7Y<�{)�/XνL���Z	�?�Q�����q��$��@�Uն�hw������6���V�ͫw�'5��7@�V��"B�4�E$Q��I#�9�/�H��r�=��9�SGV+�O���K������Ib�faFǙ8�@�aA?֍7X�*mveԲ�Y|��7j��J���h�5��Lt�_�*��O�ϥ�}a���8�2��֑�m48c��?=ĥ���>lr�ƽ �����}٢^�+����{5��>��"V�u���o�g5�=ܲ2�1�7э�\|׫YƑ��i�lըO6s`�C36b�eFQ�sHh5:�*'Y�}z��`a�~
�w<�s��p]�f��:F��m�t�Z���:7JH�˫3���vp !���cn���㉶����5�,�;��K�a���ƶ�C��y�24;\����̮4�CQ�0�ҋ	�)z�2��A�Vz�1�+/�D���]h\@󆁄�����oa|��х�����U��P:}�����Y�ު���;�c�F�&\�"G`*�q����F�XH^�x�ӡ������B�`�����A����+<,��O`�N����@aNg���@q@�m�ub#�'K�$N©���P$)��2g��ߜ���)FJK�WC����7�;�H�(Ig�4&6x���]pr�A�� :��7-���#�����-���0������"��- 93��P�RbF�/�o[��X�D��_�!���|�_"g�j=�#�;� +�qH�Ol��#넓�H��ʷ�F��G�����>�!N��=���A�
Z3�'1Y�� j9fveL��Z�â��:>�[��щ�d��o�k��^Ec��g[����3��!HdRgߦ�ܕ��<�W�I�&���r��Yؔ���"�P���PU��Aj�"BG2K��0N�[_b�2A��&�������<z�I6�;�]���~ɭH�N�F�KŴZx�e�3&��G�sZs��;��R=U7���d8��ɠyN�y��&_�O�y \��v���P�O�.99����΢{�v�>�q�iv���t!	&��~�E�3(�j·ӒQ9lJa��V�f�=՚��:U�h�RAu	�ju�3��G�$>b6�FWC�p�گ f��)�����+tC�-�'����]gդtO�?j�n�� ���}R=�<UWw��y$���Sb��o(݀$V�ѥ��V>N�,�Z "�(`�������]�1��ϩ�=X�3<
I���de�h^�q}��� ^���t8��˒P�w�q�i���>6���Μ��E,���5�d�ݍ@6p���ѫ��ڑ"��>k��f�e�9���������wņ��v�x�>m^D��Ȍ�7��*�1�fL�e4��v�ϫ	_�h�M|L�9U�;�t�
h��L�L�^nr�V�o'��|;I.S��%����@���P!L��������g���!��m��e+nV4��z��A(+��鋸Pu�nO஌�)X���~��I�{�˹�!�*�Ԛ�1��M�a�q���dt����nԷ�E{	�	��8Pd�o;0#�P"v��A��pDN_E~�����\�6<Pp~LW[��,P��%�mT`��!��o<�h�x.���fU�HJ=+Y@(T?����kN��4S[TCWB#=c�7@���4X�E�kmj"��:�U���6��R��:[�Q;��'�!M)����HĜ�%C-����<��>��>ȋI)��#3������P�-�/�#�|�Ű��x
�F�8�#�{D��Y�t���Ǳҗ��Θ/�3*|/<�	r��/� Q���>�;p����&:L����\BW�>�}��fڣ)"1B:��@�Ⲋ�Q�1̞�B�@Av��)CP>��-~S�ɒ	�)T���R`�:`(�Ͷ���2�L��56�Nϛ�_6 `�	�}�`Y���I��: {ta��*h���C(�}��G�\�K/b�S���AN^pO���C�%E?�i�@� �v4�[]~?5舍�C�0c׻��j��"��=���kǪ�@ &����P&H9��Ņf܇R �t!G�0/�ިo��~>�\G��YKR��ܡ�p���ب����ٲȆ�Ob�04
�yG��GK#a���\k��4#-y|~�؝Q1��>aoocu3�������'�$ڠ���X��G��`����|��1��O%B��P�vp�o�CH�&��RX�	բ��2�OFP�?dqb�H;lo��0�<	Gsqn`o���;ǰ$(غv@����"��&�ޱ_NH�[v{A�)�c�"i"%CS�*���#q��w��q�e^�pw}ҍM8i�g����?9W�D�y�=R��4U��[�m!�ø/;��W��\��-��>�qmiD�X"SaEG@&2�#U ���Ȟ{��߅����=b��a4��^4��:K�K�Si�D:��9E�L����B�F�̪�뿘crnpg�������z�|��.?+f�ɍ	q^�B]ˎ:]�_f��
"�~@�.	1�T���!C��������S��.��jI�,��p��t�/e.�n����x�~�GA�l��f�*������]��$�4��MԵ�g�o,o#ؘ�����3��Ex��أ)%7�Ǧ�����M�T�v*qg��x�~��@�=��#q}�)���7#��s@��ݱ(���n���n��rA���}��$�7n�=M��^q@_0�I���P�`لΘ�K��h��ATU��w�\��z����Cɗ�s��V��B�18�����H��K��g�����%�-�=W�ZFt>��_&:	��Z玛;^	�%�J6a�ݿ���z)-�!rܖ��F�����\$�A�Q4�Z3Y1�l��Y-:k���3�E)R�̲^١<�q�� �i��_�$���n���er�.�4�;/oU9=��L���W���H���N�ޝX�s0�u2��L����B5�irc	�p����k����=����24�c��ᚬ)\'�U]&�?����y
y���g���}�]EP�0��|K�fz/̰ �h�Dٲ���,�-�;�sH��Sc�Y�꺙Yti�Y���HX�i+:��(2�myX�C�=��@3�����I����#��[;�XG=E��E$Nv��>fʎ�k�g�y������_�ϒR�$ �Y���N
�n���1�e;��E�Z��R�7�xb3�4;�{��]B>�P�=��j��x�����B�+ŻT�O9�̫Bi����3�.�~�SZ��1إ澷Od����"��U�#�;H]�iG�b_W�ͼ���(���@67_pf�e�)���hѲ'�H�V��#�4�G�oOP�_.V�J���ҋ��5��̓,\��$��=EkM����� � ����I�ڷ*]8K4��NmCbW�>�#;�^�QP�)����E%��lH%��(7��4M��V�3�g��s�E��,�TE�.~r��샌S>�Ň@ �[���i��_AH]u�H5�k��ʹ�U�qT�x���b.N��Xm��bF[jR`�� ���;�|~{��j5Էo@ƪ8TiكYa�������D�m������7_�����ՒM�b43���$�|�4�*����q�c��C�eY���T�"IY+�[u˶��)ۼH���ž��.]N�PS|`ρy0��b�: Ŧѫ��[����t�q��H��$�|Xы�:㢫m�o90��q8����s�8zX8
h�5O��S�Ow���
9���#9����V&��<��XH��%`�Nx=�_6F�h_�P���9|��D(z�l�Xc�T;^�����Z^p�bK�o5�_��L1�'a�>ҽ�{������r8T���=��ňZb^¸K(e�a(�Ჱ�i_�P�
(�����]��p�b��9�T�K�YSv�V�f������W��+�ʚ9� u�1\��^3k�%*��s^�%��2a�ٙ�?A�f��
��[K//��1�1�]��z��f���j|4mm7��'��X�$2M��A����(��j;�Q�&hu1�@���hݐ��s7�/�#PR����c�;F�B5�;�+csJS�-vH�3��A��̄��/�C����iE#�]9�s~��WOkzm5�v�xOJd�T��N��eY�ds+k�
Ϧ�9�Z`�9�ZF+=��P�R��0#��|6���}͇׻;
p_���`L�?�dJ���6*XH%~�-���,!4��Ƞ�����.�s��H�)�Cկ��m�bॎu����	G�����K�>��>A�������K�}��]'��n������7�
1��_�>�/X^�7��q>Q�`���X�l�<z�H��L�q7�Z^��2��!��k��$��q��w)�.�{�MӖԳ܎U��GI���/����P�h�'�S~���)��0*\�& =�#rt�h1Y�4`K�)+7�w����5N~E�s��L�s!v���W�c#���%�����F��s��"�W��Q>c���B8V�d(��q}�C��N;km�.���>�6fbV��vY����.?��w�M������Yڙ �5{KpZvo�>\�:&9"�� woƱY����c`'ȗ��+l�@
��p�eW�0x��] Cg:\���:��D�W�����-Z�L<���/y��]��^��P�%�H�:�G�әaJ����D��4��g}$��x�y�Ƕ�H<�Y�nErӽ0ܗ�Ro��X�(��نL?���+����r]��Q�ZG�����g�#�6q�������|���-�R?$��\q���غ�)Y�/���M�LΫ�v
�B���w�\��^�9(��B'�*�jX꫋_tF���Ǯ?|�UQdoN��b%����`C�:���T���k��uE^��!��9cl������)ha��}�{�<:"�#N'�e��U�}d�^�#Y@��iJ�����|�R��X�9GǵƱ�=��A��(%��cl՜�\Xt[�E�"m�H Vm���A�3T��NM=��ܾ/>"��ϸ�~����?4P{�����=A��8u+��CM9�����	:���$	}�����.��9�.���A1' �)�;ɰO��!{I��I�nT3�oҺ8��Cbs\z����ъ�:�=�ps��5lo3N�h@�6�[,�%�Ɣ�&:c\�@n'�1�=�@�90m��9����I�Xح�#5�[K�E'���j���5�c\������f��b�����st�]����|�ZQc�y�ƒ]��j�*=w�ص!������P߷�&����:��-K�y �ۺ���w���C�㩵�C��~��� �)�+�7?U�Y�t����6�)U�$�Hq*;��y��>~Ǵ�Xq���� 3G>N�vd']�ݐ�c�Ŵr��8���T��L�GH ���J�� ɧ�й ����F�p���w�3n~n�ѝ��U�Myd����}h�'1=�e+C�&�x�*�O�F����]����3�|�q7�kJ�6˺����	`�ߕ��(MsR��Sk���4�ǟ�I��ƅ;�d�~:�o�	�:}ˇ��尠�e��l[�I�p+Z�\�!s�2�x�$�$*�T��N��F0��>M���)�̒�z����.�X��!���ӌ�:�S�*����q݃���5��cW_[��Y�][th{r�:����$�p׌��:�C�@��$]>%��O�+�����
���<��a{�`cI��/.{�B��[}�Qr�~�p��2�@�⬾�~��HȋTe���
�f6mlI`8{8�8�N��m&����}x&%N���0�S��Tcd������M������/�A?��#�n����v|Ax��
ݭz>i{�2�ߘ5/�	p�U��W���zo�5��>rw��C,�{�x�n�S���Ȣ���M�MJ�@�j��qrQX��MU����fT����ؖ����'�ṦU*���6�99"�T�T����tC&�L����B��x��E`�D�uW�(,��ܟq���l�I��".z�F�}N��3׬�X�Ƶ~5A�b�cW:���3.߹Z�r�zL8���|�F�"qq:T�t�l�0i@���t��pB�B�yO�¬���k��ҿ��S""3��i{�02hX����� �Q9�� Z^�G��4��y�������[/�wPтB"�C�:�?��D�0�Տ���}rH�6�Ub���߆by�b!�~�Ѻ1��� �L��V=����*Ypn��Ѫ�{�s�c���ND��z�*,�.���%�C�jɿwFzw������#���Z���M�U׬���]A*c!��Z1Hu�%^�:��[���U)���Ϥ�bR����;�f�5���F��T����b�>G�QEl٧��7�5���w&���.g^�>e�X8�YMUY-J�Va�q;�c���9���j�"٭J�P�e�q�M��+�w��D�����[��:q�?�?�l�ӞO|�*��k|�_4�4��!�b,�ϵ����p��/l-Rd���X���v�l�~�"M�4aC{���>��x�L�RX����/Έ�^o,緁6G��({�3�ٟt����,�"�[�.�b��4���L�~�^�$\z�=@���&̂��c��� 4���dU��Y�3JP�u
� �BD��W7#<EE�i�5�a5k�Ag�g��Z2���A1E��3�����N��T?�_LB�5av8`:�p�ϒ�� �� ��D����.�ݮn��
����_��_O�,���"4$C��j�-M�^�)@/�Ԣ4(Nc�5���*�"���)�w�G���V��R�6>(ؚ�b=�������P~�c�s0�/(n��!G2<�&BFA�|f�Q�M�.%�#��R�b�d�$rL��H0H��=�:�ʧ��S�6@����뱦vYY�j����ɡHY$��V 7����J'9��Z�Rդ�9��ޭ�4�˹sx�A��r�Q�v��"�Z���+ǣԉ�FC��Q�~	�����Y>�R��3��B�����:S�]�^�|O��g��.2V��[2�����V�BȦ��OjK��  :��>���kA>�N��]I_ N�n��>@~�����T^C�k�٤�l��0Vn�o'�/�RRDG��*��J�^��2��:��w�T$�Xy�"u�������A���"Ӷ��#�%����v��DL�	���/�G��Z��D�ހ�Of��Sw��U�z�	�o�3pJy@lLw`�cvLB�c�A�&Z�W�3��&��L�H�5Y�!��I��T�zC$H]�l�;�J��%�Βly�t�v�b�N���l'���q�m�1w˰J�!�Y���o��^<q=��T��k|��ZO��*��N �� >o[�V�}�h ���=p�&��~����ZN`���ㅓV�_S�u��}V�N�򕍸���p�n���5�e��E�t��H�;@,KB��*FypN�_����3���]�!Mq���sXx�^]�k���E���L?��0�σ��X��8�k=c�kj�����=��(���������Vf�k���>�O�Ƣ��Vj^�ڿ �|m���e�-����@����tN�i�T�����R���x�VI&��Jb����Ƅ���2���D:�)l]��H"�_�����b\���?8��i�K���-&�jE�<�*�|e�!Gt����"T���^�Rɰ��㣝�}�̰�c_�йg��H�(��ֳ���^9�%��Ld��VeA�.��������F�s�;�[\*�*V*��i��vI[�o���4��>�\D%���%ܕ�3��;��VS��俄ݳ��M�kAU%��46(�W�`�iԓ�N�l�/���4�
C�`���m<��X�֑�^��#*�?6�\U&�=E�
bċp!q��Z��8R�cd6�
���XQ����3��[����I�X���eHgs��h��I�#}�2��|;GN�(�e�H�eh����Bİa�TAG�6�$����X]�qߟ�/c�!ȃ��e7_�5q�����6WRF�y�X���$K)�RjZ�֯:eѡ�6�go��y��¼�vְ�*��^���(7k�mr��QX8ᘴ����e�e���ܹ�uW���m��2�>�������d��H(|)��J��mЄVS<()����q��&v��.�BM-$=I�3��.�ֺ�©��6�k���Ȝ��^�m^=ɈA ���vjy���U껱qP�eOIC[�-�K[��P��y@AU���n%gv���v=ȣn�}8�y>�E1�EaK,�3*���L�2�>��VN:8T,n�'==ί���������c[
��O��8ŏq��k��}�p���6m���i�~D�JMXT�Eپ�&'y��u�����k�`n�~�z+j��#�>�#!�9���,��1�x|p����������R��G&%K����2P�MO�2�7m( �~�A����@���>��F;���2���ַX�*M����0�h9-;�7C��^�6 ��n���[=P�~/�;Ѓp��t������n�A�Ym]����#Ǽ�aE9=>P��#�UN�lʣ���5���^H�b�:ZH�.�@b/Ya����XA���=@�
���ŀ�km�>�>1Pn�1� A��E��(�K`�u�� e��ԩ�@�P�ֲaD����+��������6�q�R�ʥ3)��+��{�� ^2ߥ��N�o�g�Ъ�6o'%)���ܷ��+�5-�|�j=4��{��O�/t~����r>����k7����!,�,}��\3�yc�����B���BP���3�h��Ս2��1\�l;w}�����Z�Bb��D,�������z��m֕�Q
*�4��ǽ�4��ђ׈G-Â�c4F�|�TA�[��C�����X�]����ǎ�&ZY+��yg�۾n�"x�tj�H�W弳t��-�$�Z�
��9@R��և�x� �Z����v�b�˿��Q�sS�O���b�rZӗ�JVߚm��k�:���ۍ���Yʈq�Qe�t����?	,g@��q��&l	�q���8a���'=)q��T.����zJ7j�V���IP�K���b3ĝ��o�{Hƴ���W}��iG���(~8��lb���E�R�t
o-T����N����KW�Pqp���ZG�=�nd;o��0�d��k��J�[	2"����5A�� K�B�k{�D�C�Jp��#.�������4�-��ˣ=���OPcc-�|����Go���{���𘉔9�����4����?�A�%��D�ť���bK��-G-
��4�?��p��G�$o,Fx$p�ca���ɖ+#�����Q�I��G
f		��i�㶖)�gG�_��M�:5�����oC$%�0@�̇��v1|�z��U�0���uN�\U����Ц4�f�3@O}X��eB����I,-4�����L��u�{��$r�#�
S�P����{��^iT1m��:�PsS1�Tǉ������m�P	){�Gko܆���K.���H��w`V2bt�]#�{���e/6�8���'O��i.7�Q�w3���b��7e����,+�1�}�']�%��@0y�O�?,�ʞEf�~޻��EL����oQ���<�x'�wd�,n�A����ҿ�;-g4���\�.X2������C�a�;�2�)���|$7_Հ�,��E!���w��e�#C��g;��S��h�e�R�<
��@N�"��͟����RiÞ������w9hƴױ=�y ���L��8�\�J���L���9����ҮO�w⊐�m�S3G�+���e.�����!1{��Aj`����������oM�=R���hٯ_���I4���x[�g�c��H�#��gg����O\JW����?��%�op佹�?�#"�Jv&8m�T*}�_Y��!f-���u>�A�3O� �Be��ݗs
�� �>7^Lb��%v��6rU�b�ک%?Fh���-�yas���9Pv\+����:��Ax�=@#��z5U�yv�`�I�V?`ɉ��:�;[^����Ӑl:���Nu�����(d��^�P�����\���,H��$��AB��
�����������$�޵���3Л=ry��}�Xc��x}u@)?�1�����n�(��C�m��U[�/U��v辳k��-;��*�LB:��n�M�kt���k�E�x��h2/\�ze��C�Y3X�A�D��*���,�O�V!fɞ7� �������܇���V@��f�u�H�)(�w���ﻄ�G*]�ջǰzC�I�N���Vs���Nq��MQ'�dI)�V�a���kf�/�u@Y�ªBE A��]W�./��7d]��Dj���o�%��oEy�9��mS E��KGg���(�������?�Û�����v9��@O!�\�8���L������o�5�P�6$�ME�8����4�$�J{��w:���i�GY���a��M�Ï���UR,݋���Y��PN甂���`=m ���6���VI�S����[1��آguR��<�s�e���aTv1E��O��V�7��(���j��Nc	�@��D��hm�H���[B��b�YLS0qM�˻p�@�=6N�}�D7��~]BϤ4�Z��<��v���i�Rd�5�@��.뤩������O ��LS����ՔDM�w �k����o�f)C�����3*v��Zo+1��$��HF�V�j3U-���a�g�!6��|a*x9y�@�:� -ĴPP�1���Zi��E:TeI�E�
���5�_�w8��^��Q�:�c=��X���5wH)�����é��(�7ںR?9�4��	eǁ����ͦk�Y��4	̗���3CDM�Ho��A�-;���z́
m����H�-.^�%̓����7��v���� \ꁙN�TD��`���e$\�!���.C��;��I�J\��Pz��=Bh��L�ɼ��E�%鶤��h�}�"��E7Vr=�����!�d:�m������1�����2%d�l�uT�X�
7���ӺY��	���A�����>�R���C=��*�]�Gk4wux҉=���e�1�>�2^������O��B��{5���I������%�,�&���'�)���5����n��Jgߞ��,�e���|����f�E�.6�v��Tq9�l��nv �<��*#�b�M��T�/u���D�R l\vF�c>ҽ~ ���4C?ڛ<�CK�?�/�� �OJ�څ`��s��sb��%�����n�:`�?���1rL	�$�pD��⎵D�7e�+oyO�v8�.L,鈤�V�L�T�d��}Bߐ�[oK:#�j���ݸ����g�$ptӜ�~%� 9��X�ZM�4{���ZI`�0� �%� ��{�����޺)t���s6b*�-�[�@k�f��w�Ɲ��h�]yT+5W��I�g[ �Ʈ���D����F��=m#���ss{���P�z����� 3��;3sw��- ��c��ȿ��ชP;��cZ��/*5!�����n�H�������E!��G�x$�.�#v˭�V��6�ܔ��}jj��f�}X����+ۇ�8W��o��H�jt��
m&�[��y~Gk��Q�c��	�*����o~��^�/���9��׾x�|ű�5�Ɉ�'�r��YU��#�	��S�����>>�t���xbUo����\|��1���D�s;j����U�]Ĵ��m�\��E6��'Lr���ds�A��0��!É��j��g>���Z� ��y*��vH���_��/�ySE8X��ޡj�Z�,�y_�_�l2%��?J�Iv<�O!z��ʁ8<�COؓ�2�w=�2��B��"ra�D]8o<��M��E��+�z����&{7${�`��dt�#k�m+�B����i�1b�;�1`}�v���x:�J��~�h�pk�i��${�;�fV)\��yඇIL���#��v�o�A�bb�2M�^t���M-�"	?���!d&�{�*C|�`��6"��9� �|�9��U,�3�[�5A�Q��&}D��$���"��\�P��-	c�k@E�Ӛ�%?��D�v�@0����l�rƧ��bC׵��@��%n`�@���������؆�������c���Ţ�<Y$�'���0<�s��I���l�BOg��N� ���/�r}��Ș֊��7TyZ�W�a�jU��A0�fn%��b�ENȺ,�Lt;g�ڔ��ׁO^g��٠n��&%ա
7��ؤ�p�8��U�wt!/�űN/S{x���*�=�#ՠ���]A���}n�P/4�>�q����[���Eca��+yN� �� ��Sj7"W�M��ۡ��O<g�߼����"��_C����"<̓�W�t�K�]��|POZ�W��F7U[Zd�lyM��%W�%o��������t�t�K�$���6)P	g�]G#/p�tК���X���zp���ʙ��O�G�n�������d{�����ww
��;��e&��Q�[vG��b��z�������̭��5Qꠚ&��vB�����xS�ͯ�� ܍2*�\�F�@\ZI0j��uou�{�6�L���8��V�ώ'J�4I���uJ$cva���[�J�u��]���L�鞞�6�<��&�����t�3�s:���@�����v@k���H�䴛V5a.h��?o�~ڛI�ݯ�s���v�r����tO�Hۮu �M�F�@k�ި\+Đ�2j�P�9k�6�7��2.5t���<�T�T6ż��E��A����\�E�zL�
��$6�#�M��/���e%�OmJ�p��Z������(X�Ҏ�o^�K%]O�.v[�C����6~����xXF�y���!AڢOvb{��a���7*�yL��qE�� @�`�!y�˫�*�]N�1\�Y6]5�6���z�����A��[Î�$�+AVG��9�p���'>��R���&�S\�'ٰyk�c	lM��>�ā���D],�����	=����u��S�	 �v�G��~=[~�ë� !�E^H���.y!�8�I�d��I�%�Vn�9�������0a�Z�ȝv�!s��Ҳ��#�0� B�r��_�0�W:�� ����s�G��"�vZ��O_�Xjeۏf����1P��Ok�C\��н�Ĉ�o8*i��D�0����d�~�n�a�In-	y>`��Qb�߀��%�5r�ӣȽNO�B
�倀�E޻v[/���B�r�PǄ����Y1%m��mv�Ԛ*mB�F�'��+a�f��m6Z�=�ԩ�AKjM9��n��`N1�+��('2n�3��$	NVb�����{�h�*j,�B���ʽ�\T�N%&Z���R�o&0'2���2�i��P�u�g-₠�U��!�������&n�@/��Q��~� �e!���#'1w���tډr�
�K8Yh���o1)��Ibɸ�B���Y �E��+<���aQ0�9�2֑�@�����r�Q���թ�O�E]��� ^��A����I7� ��S�<k�����4���'X���ѲE˭��~Nd�|��/bh��tȎh��{oڵNܟ�%��@/v^8eޱ2I���$�����3����;�(�N����aL�����՜.�ꋡY��b�&!�f�:�\Z����W��΂�I���vCT�F��y����7u�Q=Wnk�P�]�{E_����%�"E_�;�����Dvd�� ',�z�@c��<ٮj��lx����H����������#&w�'`*����3�m��a^B퀺|n�?q��j�M_k�[W3��Nk�+8���!�F���[�t�Pl�Kt5��͝2��V�)���Qp1w�D/3�B{r��I�Y�_��h��+��ޛ�>G}��ae��+�oL#��㛫� ��Ǣ�Y�@t^��D�^�2�?�$xvQo���W����K�o����B��{?�(�ċ�G�"q3�si�� �7s�16�T�~%�:N��3fw�:��_�� �2���G�rHU���v�.�%7߃��Jt�����`.��QQ�Q�J�U����M}�ɨT?��Q��L$�����B�s�5�zI�nK5j3Fs ǂ��=j4�y�"�
~J�J&� �>,:#@�I��`)��W�^�\l̔<��bb*�Gqt���3�];-G'��&Mdy�L�~
�琢뷯� A+_NKo�O���=�B7�5�F<�mA^#^c��TI�*�?���4i��n�ƞNe��T^�#�F ��l��4fT�Fn���p���-R7�l�H�j=��C�$̏4[]��<[����P�X���y/X�4�
�G�VnD�a�����q����8>"ʮ��8�,�+�G��4�%�7 ���0����_K}R
��Ͽ�!��4���#�|�-��=6c��~����s��lL���8 HB���	�Q��o�h��-A�j�,�P�Z�z�'3O�Y����=jD��Z�\�O�'�Q��Lfd�ZX�P�ޱv�(��!�&U�4 ��˓d���#V4d٭eA#k�7�%���T(P-e�d�,�F]���x�NA�ѐ�'���/ކXy���Jr<���%G�j#�a]��Iא�9^<�M�w##����P?�].Œ%af�>�U�_
�8ޖ���[����f�S��ANe���#�m?�R��7H�"6s�Hx�7�1s,Q�ܾ�����j͟��B�_u�=�&�9�x����ąN�7��r2D���7}9�J�9Y?倥�sX��J/9m/ˢg������ԏ���d.yИ�Ɠ��tf���'dֶ4���^R����Πi���$�����{������G_=�p�=�M��� [A Қ�C���%7���M��`t8�aK�b�p_���eaMK��l+��|����`�2�HrS�♵�pt�0 a{����9|kS�{ݥ�^�Oiy�
�M��7�J����U�N�]	e`��'&�A_��{q��1.Z'$0�e�l�*An��J2x�R��C���^O�
W̬��<����/=���r�W�x�'L�7/�'�$iW�B�׺����ӓ���ɐW6-�LP���s��J��*�,u�U�=��1���~h���P;?����ߏ��G�#��4ܺ��a�����Q�b�F�U@Q�P!�q�N���E�r�E٘+����GY�b�r)��=�H`Y�w[7�ϴv?�v�۷E��%z��i찋@��ߝ�����Ȧr��
�^�'˺UA�-V�ZQ�[̤�Pv2������!�L��3�Ǡ"/�q��-�_m�x�6_�d��\l6�8{���j�z���լLj��3U-�#�}ź�a��Q�G?���LQ���j��}+IO͢�����7�����8�Q,G�mo��-�bc9�*W�h�� �G�2~�)ϱ��\���x��c9ĝ\?��c�vѵ�:E����N��#����	�s����f��o��|����\�7i<X�H~�eD������ �r&c}N2l}5����(y��~%F<IV`�@j{��6�����r�U�c㲇������mP��o�r$��$��L=��Ƃqk��������JJ]�-�+��r`K�H��z}fX��m�k�g�b�#r`z2`�\�i[��=ˤ����12	*qņ�_[�%�`[~χ�8���hb�-fo�̵1O,�9C`z�V8��&�F�!���t<F@�w�
U���ԇ�����aLCuNV�Cbq�iF̔����9���c�S���~'m�C>�\�{"IG��Z�HZ��Pb���I':mf��o�V�BȪ�յ�q:i�f����a�p��VqQ�	�|�4J��]��g"��ӱ�-�<IıI�z=�S{�iAʅS���Zί<Z�Fd￿��V�7k�oٺɬ�̀�y-����CL�������-�4�� ��C2���]Z	l��9�T�޶	K����4m��%�.�Q�QkV-.�<3�js$#6�d�	�wi?1���d8A��ʨ�d�aK̛
����cō��+�I��1����iY��k[c��b��v׋�+=�C$������֭r]�] c|��&gi���J@[�8{�N/w�Q��$�-�4��W�tS�2�H-�³g����|]�K9���z��I�Y�Y�eO��@�W���mH��PY�ѩZ����iv�h*�d["��p���3ի9����~zO�W �ZI�w�V���ڻ�V �"W�	HٳG���o���PXu�{NѾR/����g���a�nM��h�L_�����?���^�89܍�E�iT�,�ӂ�y~PkF:����7�@��u��z���^P0?b�'��p�K�}d$���Ė�qM+II�B:�5%t!�H6�FF䂁\�D������[l&��2�di���>H�[35��G3�^���~��u,oky�O�Dپ���K;��֘�e����
��H���R�t#��Ն5�o���:V�=��`6��s��k���T�?l�������wIp)�a�t��@�q +h^ŴI���
=	@��+�G�&Y�!�߉�����C�`ŜP��q+��ALfߐU|y�"@n��l�F<�`,��0�|�b<3ƅ�R� )b��-X�5]��ߢ���ń������@�_�y�f?`yK�A�Jy2a�>���s�:B���r�� 7ϊ�7��[%���Ʈ���<�އ#�ف�?�f�9 7�ʨ;�"�6W㊿@S��/�'u"g����ddU���q��-F�k�Hy��\[H��Q1x=�hU[��j�q>������>�L��:8�h~N�KԊ�CW��(�!	I{K���t<I�k'|vBh�i��]<b�o$G "	'��V4Y ��9�k8����.6�Re�r^|w ԧ�k�	Mde�OI4������	�3$�t���R��P�Ú3�j��C .�Ҝ�f��I��D��?��K����-	5�{ʧ��#6&^�]�ź7b߄EB��)��)�w�� ��!�����ҳ�*:�����S8����3�Q����S��-�`J��Ie�g��Z�$�|y��LdfU}u6��Dr����|���ί$i��s~I��A�]�쏹�OuoA'���vZC�\M$_]0��h�^���ל}�y6��W���1r<�,8��� g�!R�6�Q�c:F6�a����J��"x��M�Vя9�|N<���{a�J��3���%c�1�r�W�p�W��S�����	����Z��d��v�2 �~q�����VG,�p�����i<���ۊ��n�������jm��`#��7�O�`+�L�ěI��'/���P�$2�����xKή��A�3�}��ңn*b��%aKF��6���]ɯ~�H���]ڴe%��o�3T�r���r�����c��&[k��0���i���\��9�:у����n��=��҅F�J~�	�@Dzy�F��ľ�t�{4��Z:E����6��u�Zo-]A��2P��y4c�� ���[;����3�`3�I�J� �*	BL�vi�,]L�9M��W�A���ë"�L4�;�HK��&C�lJ�v6��Z�1�]`>4V2��<Z�>�לw��ᘅg�(<s	;k��e����V���,�Et���8N0�u�Aj;T����~�����Q'=�,�Ϲ0�#���l��'nAI?�l�G��U�B$����PO
�kN�~��7���N_�~��׺"���=Ҏ��5����(�`���f�
j��6$�E{���ɫʇ�U.S��_�J%��ۓ_PG{0n"�`O�����Ћ��vha���A��e��i|F�q��듽Cd��yfz�݅@�c��%�>|$	��@�C� ˉf���0CTQ��Pz#�Ɨ���,��q���dSI��}��{���p ]�V�����,J���beK��X���C|�����cE>+��IB�ԝC��qM露S�6GP�N��m��m��.�K�2R%[�y��;���f,���I��Q�&�2��f$��;ä��p��N'���X+y2�%��K�p��z�����X����5.����Vau�>�f���#��� 6-4��t\o��w���.XZ�lA}p�al��M3'��֎��N�+�k5�`�=5��iJ!9u#y�H�I��W�;��J'9�
��%F}�Ã1�ܙO�#X� ?¾�8$c=�=���-1�����x*�摸~��Nl�0���ӊ�n.57�|C�S���ȹVu�Ձy�	���1�&V��n4��c�E㟑b5
h����1*�ה�J94���3%�w@^����,D/9T�f�R%�d�eM�Ţ��t��0�HN/2̸nFe~"S!�In��E͆�����c�ڹp��*R��̚�+���2�O��Ay��~����ה�g�m�t���T2����g.	�h�Ӊ�_$��z(�w4�oo���tlRMx+�򜪏c��t���(9�+x�J`�UV�,��S�Lt���箙L��M!װ��d�i���Uh�}�4:������V5��N�,ZXI�����#N�_�	�=,d��7;��Y��ׇ�5���(���F�����r�q���^��kV����g@�o��o���N �����_�=��d|h:k���l����#XOVѽ�%x=�Ӿ�<rE���K��� �}.ҿ�F�� ��h�����:T�w2ޱ�9g`��(��GŪ�Z���9����<\��('Py�m]��#`�n �N]��B�#�ސ=rZt��9DKn\�1� �8j����5VW��̝��V�5 (���M;�x|�\ծD�!^�2D�0;�F��kЃ��w�'��>wn�`�](�vy���y{���\�ى�������-ۍ�>֏����q�#�/ЅD�M�} S���l:!�������G�qWDw����+���ӈw��(��z[2�d�ɥ-Ku��2�Pm0,*�4q�N&��2�Kɂb���K�)w.G�K���جɢNWR�J�����2l�2L���pqB-�-���<,�ɭ��gf�)
B�c���,^����g4�0Mma�}K�{�6v?���:��>���Qm����9mr�"�x0D�E�Z�^qSu.�5���i��7{'6���I��}�%���~7�ַ�ߐW�����k�!ö� ������U���P\a-�{�ң�K��$N@ 2�|��=����h)�ص�d����W{#�yo$ʅ�w8�H��y^[��E�|׾�����Q���ÔnÐ�7,X�ɩ	�Q�i2�	Mq<��u(���<x�%�AA2���-�$�!u��~�}�jh�a-z�η:�ާ"PQ�`я{�#u�����}���[W��Uh� ×��C�j�
0��r��o,Q�׌�a����wLt�M��>���L�y�G%^w	|k�?5������^���\9@~9x��N��N7�;�Mv]Rƀ���w*��dk�����G緥���P�1��Db�(�M����f���T�2��	�k��J1&)��(���z:,�Zu-**k�"k�D,���[��9��u�'�&����Aݕ��)4m���0�+�u��{���6U�E	26T�\�|�O c�8=ֈLP35�܊�%{����w�Qw��綹{�LY�G07b
�9!Ƣ�0Z���Mbu�w�����@���)�S6���3�Ƹ7��p�lE���8��;8��?"
���#T/O����eX��K <F\DusJ[HYW��1�N�I�D<zB�v�#LB�E�Ī�����9���j�A����5�)7g������W3p�+�:2�oZ���<��g����\�.��S�䉈~�����s�`��o.n�]I��T�X�_ػ���̴�`����A�$������D1Y��"9���ޝ�y<�|�6���6n}����3[QP��e���ב����V��-�������!D��y�%���T#�^N�~��w���n�<3ހq���[Ee�M@o&�/IO-��HI��f|�ɻ �ô 5�`[_�D"	�>C��#�O�ö���5Y�]�ArŰd����
������r�Gމ�_�ٿ���m��YL�@s�N���+���kp��y��K��ؤ^s�_KRM>������*, 6 ��/��`�*�m��6��Y�RS�c�E�o���p�;�K��ec�mb�=�<nqn�$�6*A�}��܍|U��M-GZ��Xz|�.�k�������f�hV��x��z�`�m
Vv�(uP����x��~�7�����iy�ܕ;6n6T��8���[��N߁}{��9g�f;�v�).A1����'��R:s�7�\o4fį�U�7�m�e���Wt���m�䨔�+	�Φ�f�$��~������H�ds9HPfNhte����親�%��hn(���C�N�[���R�9�.�88��)3��d��&���lA?�v��H牳}�J�%�����v�UK���Ş+kgSz������`��bD�ms��m�a3���s�h9GF%��%l7m4��dyޑd�rY�$ӭ���׬��[\k�OU�$?�����!m��\�3�Q5�c�4-��^Cc�P��:���V�gef+�\��;�w�r��Ek
W+��.gS^B��3%���E�!�wJ�aXEF@zp_�Pw��b�|!�4Xm�r��2l,$�+1��kۇ�c���ҷ=��oʤJEm�9���q����R���2��~:���0X��Z�������.!�4�cjNߨ�ZbU�:�� ���@�����T�Y�,/���gn��I�l��Z�CU��gP��T��O�\fs�uaѸ�8��8��Yp������(5��}rs�8`�8�>��I)ﺻ�����*�8�rp�Jwr`�CR ����T+�ƵWX�=ڄ3���i�֏�R��DB�Vd�)ވ���������-xt�w�1��F>�O�NQl�\�TD�f-���Uy�4��v�1�W8L�փ8d���[��(�jz):i��)��	�3�P�Ҳ����Õ�M?�$�?�OL��j<�m�1_{�q�="+�
����D;)�n�b���J�����E�B���
��S�(�l_�ٱRڀa[%��#T\��,}o�ήT�I�nh�%�W�,4�Y�;�|G��^1��u����rN%j6j�L_����>�G��=2���)pqB|%��?\����Ec�h�D7�%�w[w�ʍ�y^�b�R��S��L\`�E�������0R/��)'�Y
ʺ�k�*��Lx��pM�:	��p�Г���4z����L����|�_�ٷ�M�������^����e�=�r�,�YRHW�����dYP~}~uİǍ�P���D��H�i����#��̧2���Dzֱ���(�S-�Ck`�tE���p������F:���9�E*�w����Q����l,�dx����B��l��ӟ���Վ��,�hi(#8���B���0�luSc��7$�u|�*&�Sŗ�_�����u�����+)|����-6v��H7��\D߽Vr.F7y����J��n���) ���2��j}w��?�%����~wwK�W�QQ{/0�h�o���N[�eI���r��{<�t΍Z�Cs�����QW��3�x�@4F��ҭ��R��<2<+	_F� �V�n����I+hB�����^�?�}��Џ��{T�"� �ȳ�c����j������x��3��Y�5�߈�!�իG�z��<�UPz��m$U):L䁭�*]�K����Y�hQD���U�N-�4z"�Y=љ̓�=�Z�(p�O����2�1�bſ��Ӂ./�ͣ�b�_�*�������tO��^����D�.�-���Cv�#�>�¼4Z�u���?`��Z�"�����p��KS���,5�܏9�D�9��_����Q6�ccr�P��,�����+x�w��ֶ��EC������}�?��7p�F�WW����(��P]��}nj�&�_�m ����l����	��=��qn��p@5�O�)ӴZa��|{���T���?K��6	�M�F�s69���磤�n�ϭ5<q���3�^)|�D�TC�]����d�,E�Uu���M�b����u�͙��^�'��:��`$�>�A�O�<��Z���e�ՎS�Q2 .��`T��� 8����2md	���b������c2i�i3'6�&�o<�[2��0��xg�L�1�O��S�ׇ֭Z˹� );.[���,�1ˍ'=�kNM�:�o�mں��\�b������<Nv`��ˣ�z3��Y���>K���SK�B<��{�ӷ
T�DJza+n���y�2�Z����κ�p��Сq�N}�PY��(����(�0��])��o�HҤ��x�b 8�`�� |�|�S����T�� gs�B�iZA��n�y�6rŇ�_�o���b!=)|�s��(�$�������Rp���sn�r�ֶ��(W�C,;N�'U=�DA�n�]�R}�F(w-�Xܴ�]@�V?��3Z{ɯ�|( �f/_�i<k��eLMh�@��w�N��~qoh?��0��i��r ;%��L�x�>�1��E_�D�̼��X�A������=u�L�w fӥD��쐔���?	�M}+�H}���v�'	�M%ȸ�V������M�ゃ���ل���z�)�A�x�رuT�:�Q�5s�O��k�^�$d}�C�ECV�M6'Qi%�*aǗ�8:��&��sY��	�ax�9�u�k41���B��h��������a�D��Xb�5QZ+�K�m���DG�A5�Z�29�,H-spH�?�s&#VT@�na���C�_��������2���S@/UP"A���A��-Y�+S��E������k��2XHM9�~"�wrǲT���|W9;X��^��i��/���#�G׌�!��7���*���}��x�w4�v��P{�����r~���8�������o�"��Ay����XNle���sb���r��\s'�%��1x$r��P���;&�^�;����,
xE��ᦪ���`��M��m�3+���Q��g�t��=���ͪ�v��{Y�CG0xO����(���Ӄm+��#<A���p1��7`�|��fˈ��C�~<���v5�$��5)힏$ܱL>����6[��Z��x�N��㳣�J�[�y��[Jq' �v5h�r���I��kF��J�Dݹ�Yȳ��s���w#L��,Nhz�����6x���I�\�yQ���4M5ͬ��+�z���k�V��#i8��[0 �a;,�޼�4��ΈmȪjx{9���Hps�=q�NlCc��[ӗ����>a�,��ZȌ�=��k�O��1зx���B5�$�dP$�R�/ f�b��X[l��^Ј���7u�n��l#�T�Y�m�.F���Ar��\̅vĪ�����Ν�|���q�0����rm�R��� ����c� ��_��)��pq"�����9�|l�g2aD��#~�����.�f�L'ӝ��G_�eMB�U��y����"�����ń�ݥ��xr����Bޓ���\��A���'P��:���$6@���I>��Fl\hQE�71
���|��n&�|�:�J���94��=�b�����z3�#��I�̈́aAo��]?��������������A6��Z�i��V@��9��z�&�΀�*�p ��&5�$�=���'��^�GA���5�S3xG�R�������#?V�7<hP�F^g�}�)L|�Q`�-�0$���-l>��h��<�g�N�T��ϳ�QК5o��Ԓ?zP��&��9����DTA�׌��Ͽ�m2p@ư���µw��f
!�3�>1�r�f֔���B�o��l,&�p%Q������u��U�P�Y���NS�.�-�����t��V��؊z> ne�f	r?�a�|���3|�3���r��D=����V	����5�ڮ�a���*:��[�VP�8{�x����W♍���B��.p�v��3��+��L�ة���UљBz���T��"�"�L��w��[]�F]=FD<�W3��2ΗV��9Kef9o/bCu&69LF���iQ��EϱM.]��AP��/��0�E�c���=���K$�� V�B���>3�/b��1����&?Χ�i��x��WTaE�}c��|zv�")��z�ĵ�Ǯ5� �
�,Ux�'��]��J��d��>�����H�8�~�l#�Q.�`�Z�)B'e���E�C�?G�/���E�k�F��Z�>��"pn��O�R8"��r���F�����,��k/m4K�"���7k�]�P�o�A_�mO�g�n�M�bα�_kRs���ȼ9�A��+J�?/��~r@��gJ�Ge�Q��ҫ������U3q@�g���s_𢍚n�v�{_�x@><=|�]���lu�+�c�'�K*�Ü4��ָ�B�]�r88;Љ��芏J:^'�XX�����S��$���1���=~7X���ȝwYA�k�B��f��qC�-�����Ը�Kl�a���.��%������&��T�Չ�����4���J��JWJ�����Jv�svĠ�oD��Ѥ��m��䌾(�� Wc����1��!(�#On	�0vVj�ebm�D�G,�x���c���R�����<��"tM� ��ũz�5�1:��Kz}�O�fVW�����Ǚ93?��@pN^��,�Sv���F	v�}0v�H��#�W�#`�ZâOʈ���|��w�ɻV�ϡ�����ǆ��Z]x�)ƪ�I�
��a��oX�ql��3?�~�8(�A�X��|��u<���5�*���M�]g�қOE9�n�ꗗ�>s<wB��X�E)e�V 7xс��iGn��s �s�Ƣa*:4vWZ�qt-���V8��QR _Y�Ϟ��~���˅y���VFJ�Ć�ՠo&��\���:�g�m	#�ʏ�:hE��g��[()��#�`�`:��1�_�[�=��+�Ʉ6ڬ��x�{�����4 �7��3�Կd��'xE}[���i���/z��s��aP�j7�l�n�e}c�͹�/���ٸ��W�60���
�0O�:p{��m% W�������>N��nf�DU@"���A[�G!@�t,찱J��H����\����B ��n�x���Y��1�j��u^(�+���Z����/���D�@6\^�����E=:J�63�;��$D#$��'����5A�����"���� �`hQ������m��Vl�����>���d���1H]�>�!S�Y���%�mF��4�G;D���I����ɽʔ����ل�#�]��AO�%�x��|c%���WÞ=�R���O��q�.;Q�` �
�*5���#~�Y��V9�t�����a+IM<Mt�8�bR�s���s��~N��ݖ��ڂ�g
���"�u$�^�_��C �)�w�� ���:``w$x�	��ۇa���`�xPCRS�L��%���t�ڽc�H�����"~�~��J�@?.nLRY\���{��W%V�5�h	�n9�0�%������u	%qtz8��1�ȌhuO=Y�D�0��_���g(�?B�k��fK����J2���F=̺?s(O�͠��i�}<�괅�'L�`	��rzJ����x�(���n�d�1&	��w�t������GF��w�!�$��18v�v�61(���_r����I ���Гz�������bZYs�A����6��Eo�,�)��z4�Ħ`>q��������d���H�a$D ������򢿣_dv��9�Y�w��ra����ɪ�|?N��o�D�~�.ǳ�nH^��,���Ȟc���nJ�Sh/�R8�zM@�I\�}���,hD�_kf{ET礅s� Q�n �Ƹ�t��dZ�0gS@>r�n�K'�.�u�eH�w��
a���꾜wpfx�x��J :le��	1qk�I�"��A�D��i�w���۸�RYff�������l�&_�Z�Y�,�Z�D�M�1^�M1��8m�_Y1[A��:R�+,zM�9�	
j��^K�W�	���@��_!�"��~�{�6	�\s�0m�ʫu����|�kVu^plg9�C��;<��ɰY�7n=+)G:�L0��۫lL���mT�)����rH
F<�r%o�p��wp�"���n�&N:Y)4Iڜ|⨤H�W��b�.c0��N�8�B��(�A�Gk2ZjV��	q��N��9O-�%�Ϳ� ,�٦X�ߊ�7j���P��Qz�3�����yr�
�TȈ��#�f�Y�$��)!Z�a���O�OR~�_p�WΑڷ8g��,9�������؁�t�.V
����8�k�gN��
|~r��:S�����(�Ʋͷ'D�f~��w�	�ψ�-m8-j����'C�+�Y�Vay�w�����@����D����
���L���P�;�X�%�x��]^���~���Wz[�
��Zo�|�a��tMa�*�.�4�Y3Z9�zC�:^3xxyk���6�d��dm	�Xg�nbMfr���RBԙu������?6QV�w��Q+�'~���!�*y�'t����j�pv�pL�[������8 ��s�p�s�i4Y�Xo��rE��7�E�e��aq��R�p�� "#s�8*�JQ��A9�F���I�Ə����e���bnIk�,8�y�#��Y��\�8B�c�� �7�6c��h+�zX�O";�.�*�qŢ����;N�r K��uyӰ֙$#����a��Џ@Eo��4x�Yl��U� 2��c-fu����r���(*S�� �Vm�։co�]�dP%>L�WP���f,;��������=S�����޼��a������OA�`'�T��:i"�2�D��ȸMnRl��몗�B�M@�?�``-� �O��D���g���� E�d;����v.��	@��n���I*�b0f}�H���+�� �gio�I�߼	LQ�R��ܟF_�`�d�Xo[CBv�+�	%�.qn��"@c�[3��bn����2�क2D�WACǄ@��dω����.�aQ�|���Q���o�rb�u�<����Q�i��G� �4���6�B��^wÕ*�g*���z?�b{J�p��b���]�3B|�?��M���4�\�Mr����Å��������D����P�EV������jm-)5�����nK�|�Y�� uw�����j�[��3��t�Y{���g�No��쵦4RPʌ�L�rK'�r�"�먬�|�.�n��n+�7�����Ξ�#6;à��bX��o��\�yO��2������2���W�@���޼�=.��P�0T�%"�%��?kL�c��r�"���!N9>n+�g���mY�wJ���.�˸�I�:����aM��0�=CR�Gm����̼�ߘF9�r�P��<��&6���]%xL�8)[A{ S����H�S�Q?tư��zG��"�9B�_�����r>� D[%��c`+�o���I���<4�6ؤM*i})ە�̙���w�=����:�0D;��؊�s���O\�%� 3�����{.aT�Fe��O��}δ&�6D�OO���3��H(�m�U
��#f6�F%�/��������s��>��CP�_��M��u�7H0p�ۀ&GP*U��H`>Q��^��Bc�Q�6�F�AKR07z�D��]�!�%p��]���ӣ�=C�����Sx�K�;��:��C[�bܖ����t�S�.�wq��]*�L����r�:�e�3�s�0�����f���Nmp�b�ǅ�:9:	.��H��C��p�?L��x]^�˃�BA�E�ﹲ#5i�$�$
�V�3��އ9���C,Ro�GQ%j4AozE��e#�� ")��~V�j�?�#�'Ԫ��R�[�cl��|��v�o;lջV���{��w��|/l(��8��w3���(Sjf�.ݜ(�?f#�#U�]���
�Y绝^�=`|���
(^�]�rp��G���g̤�' �ap���U�,���9�[����uu��:��hj��2�搧:ďNV���}-�U�9��~�	`�
�-�͗�\�I���q`�!�90ḵ7%����?֎!��i��L.QĲi��5c��ּ��Is;��fy#vCF��ac���.{�B������.1 H�9�&*/�J��%A��J*@xT�D�ٻ�a�P��h	��Q���
Ʌh��Ŷ�n�CA�z!�	��=Rs�h��l�_i &���EM�����W�<�G��n|v��(�A�;�r盩��^A��Mt�j���eW<h�Z��
�֦���Q�YY�Usӌox�4q�x:��
�w4��n�k�K��%uF,m;2:�����Z����c��M[���_qS�t|���`�/���Zu\���0B�RN�YŻ��a_<o���Cuλ�J-���`9���O��%B?�q�_RQ'R�#��z���#��폗$D4�����
�E�H�P6��\ة�k����V�;y�R���Nzs��Rb��A�h��2��
���%��Q�qtãd6nV�ۦ�~�%���CL9�z<��I!�z'�A�t�����+��7���\ ��~��+ni.���'�o�l��6�� ��+艎6tP�%mSC��0��o��s�s��Z���?1V�Nج�F})R']d���3������`\ۿ/�I}gt�蝘�w�֑/@u�l�b���*��f��'R2�_��8C>�����mD{�y$2<7R���z��I��^h������gg�XT�!������E̔b8�$#�r"�hz���
n��O��/�u׮S�K^T�)zF�3Oj\��AP��2uv{�U��{[9,��E|�Y!M�-���Y�VTT��6� 6v� �g��Qy����h�O��F���O�T-q�`αuڌ�����Xh�e�^OBU9\��i���tY�Թ6nZ�;��@F�z&|�(�oΏ����S]b4��ËJ#V�F���U���� �xe@s��XŜ���st5���Dh$/,���aIyO�.H�(p��+)�.�D��j }�s7��H�/\��ӆ�	�%��=w��n���p���z����m���C�@�"��s�����2��A|���R̊�R�p(C��B[�?p�#؛�u��,qa���N�ޅS#6)M�f?�>{���2_����O���.� N�>in��E"JD��h���.,��yv6P}B�.���%�M�7�%Ÿ)��K��ǺK]�̔I����+�cL����8����?�[�n �=�-FqXWCg<G����J�Q7LdiIYk}rn���;4��0�*ݜ�K8B��P.E��i����S�6��DL����g��r'J��YC�m=tK��@/�&�m���>��6���8���7�.�,��@dnz�p�S���:�@^#u�AM�2���N����r�d�dp�C��H5b�P��,��:K��`�qq��d�5a,H�}�#s𭬣�ԅNԪ4��$�����Lݞ>��{�h;�j�:���v�y�Zt��;iN~�`*̖�cǆ�	a��H�"�����@�3���hiS+q� ��m߉��ʗ�C6��V,��Z(����ItH���D��F����P�jJF��?�ǟ���+�c5����8mL�z�� �э&%��.�c�H)j,m�<��j��$=�k侦g؝h�G Jӝ��m���_��t��b߮R(�)+�/2�J���p�a�z`"7�~;��c]%lmf�-�с�J�W6������^7�'��0/�i�I;��Z#/��-f�[7��zX���:&�S���\Ƨ�V�"5<L���9f�ݲ�a nv�ܲ�m�|�6{6Pv�*�Fh։Z2�ha/�j�23��/�c[��rZ�y���d�f�)�b�)g�܅��<�~>Wpc�D;��K�wY�2=2�E1f(��U\�������]����&����7y*0��S��j���7J-�'j��4OX ��տt.g����h�6�q�N��7�n�_�E��h�P�1�u&�M�*|��g��vCh����1��8�����3�}��Lu�b�ob�\ M�/��|vXA�|5�߹U-�b�QP���
o�].���.+�ޢa����R������'g\A�u��/�b��q�)�]�D�`9 ������{�a>��tF���|�yv�_�5�ѓĝ{�YQۀpo��#R�|���N��)�M���U�6��*��1��
KE;���ԷnYx��?�%��}}��7�͆/�ښz�B�	�IoÜ	`�+�uͧ���Ӻ�{Gn�8���ٍ�0O�]��Ζz>@*Z�v�;�I�q�L�Ц�y|ow�F�r��yJ��nL�$R~Q�s�~������+��p(�(��>|R�S.���߬�f��5[���<	i���lW�b疻$f�f����y�\ÇaQo�M�*���R�91i(�z�Z�88�_zyc���m��(�@#�'���gucU�T��~�9G��x���ƨd�ǰ.�裔���=�j}��M[!r�����������$�P�c��!�m+7@3Sx�qߗ*d� �3��BnPmw>��h��xi[kij{?�+ XT�w��ǌ0=�w~���k+W�	��0��y��Ui�� ��E�p#�пK�EW��ꙃػ��3d����g[L:!��~H�̶�y{:�~A�K���?���PD�\�"d5|Ы�eEZx���VS�LM;� �<�9�MB�������Ϛ�����9$��;� '��Y���M��Ɨ߂�����nu�g�OuIO�/���58�8��:�3�y�d��W�_����A?ڶ�a�u/֓����ұz ��.S�tg�X�2����e5`��ZtI�"T����Y��
fv�mj��5�3��N�~h������ҳ7験�VY��\�I�D$MG,P(V��l)�
�L��ݒѩ����#��)�&�RQ->���3�4��T��URT@�e�O;@nm�!������~e�a3,��H�Mvio3��8�Z;S H�����>n�(8>͠�7��f:<���%���Z��^&6�P����X�6U٧��T�����Y����(zl���9|�M$�9-n;���܌�		�Y>�;O&'�?K<�`/a�4~c���L#�ё"��uꑔ�Qm�@�`��%u5� ���ʷ{�u�ß��g��o�\�Γm���A;�"�tD�P"/��z�9�(��E��&�2;<��������>�k�p7���'���Q����p,	����pp�F;�z����׾��U�� W�|$�M\�z�z)�m=a*��!�JFP��W�Mrqi�O�C�.ݢ�$75P���ա�+B2��nS��K�#�wҩ\�[�.�H���`wM��1��v��	J��N��D�]�ba�iD��E�X��3�XR�<.�z��3V���<g�6V�hm�$j�Ǌ�Z��/wIs���5
#v���lGQ3P�F2��F��,`cσo��������ƻ�c�?���V!�,<PY�DP��xw�8k��Av�?�GfTbv�D�@ߏ��j@�naְ�r�e�);	��:G�U

�՝7\�`�/�F�����a�x��s�TX�I�V�{$2��x��!
f2'i�-2m��Db)�L.ᵏ��>0fҼ{I�ᯭ:��et:���n�t�-��8���a�9�[��_�>t�����D»fx�䶋�U�Y<p��ӯU�o�"������*�o��:h�T�A�%�	��E��ѣ��Y�GQ��W����8�'�J,�sK��b%�����+����F@�-�y�� M&�USd\��b?�J\�a�~PO�!6o6Dl�Б'�p��"b��й8�y���z۽�-E����=L����F�UiT��צ���C[b��@|'v5�ƴ9R��Ǟ���7d��bG^iF�|�;,�H95c�){�b2���+f/�*B�
��[5F6�`ł�]����¶Sɯ�'�=��:��m�P�;�-;�d�C�'JR�9����*/"bT�����܊\�j���&+�5���^C|�g�+�Tz	XZrt���X�7��䗟�
��e
��F�ư�t3c2f�!Q�~L@('��L �;:�3T~�18:�����C�#!=��	�RVl4:@o�ށtܡ�#����MH�}������A�+�PFe�`��Czh!�:�##/˲v���p?�e��`%���O�z�m¢��(����Man_�>C@uA��R�n������Ll%(򃪼i�q� d�v߂�H�?�OSp�ce7U{��G�!�. 9�(K�ߍ�뷋0��h��K�Q��!V�ф��|2���]6�PE+Q�� �Dj���%�b�
Jw84q0�ǥw����Z�O��v��AO�{!�K�[�*H$l!�J\������qh_Jv�筳�Nd�~��ݍ��t�Y��C{�\��t0�4��Fѯȳ~�ά٨l�3Hcvfbz*�&}:N��j�em�р�iޓ{D�_�*�VgJ^��t�m��XOG�����'�_�A摮�*�Y�#�Ҟ�cw��S.�W�T):P��P#q����V���	�k~�����;?�����%T��c��\��#|ς/�u�}��S�V`ur�SC��#|g��ծF�R�oW3?W�p݋ڠ&z.���Ǖ-���eQ�1z�7���ӝ�rK2of{��*����:
�G-�S�@r���[�Q7-�%���X��U�?2�aZ��lDu&�����@gR���p���� oh���S��Su�A�5J!����������k���(B+��[������WY2���oə���f��)�=�7�����.�>�������M���h[\@�8��Q�J�~ۿ�1��b���y<��,!ðK�ghh�8���Z+���w�w\*U���E�	 ��sˏ��>�k�l��E,�
���+~��V�����CPA�{� 䌽�L�)[�8�	 �kˢR-ht#)�ۺ��h�ȢN6z�����4%^^�+���kj�������g��
h&����B�j4܋�v�����/o(�=C )b�T=즸}��ԡ��6��b�A�J^`��$5�<��j��r3P���f;Qf���IO=��ڃ~j(��c0�<�z��u!Q�F{N�oz0��Gᱫ�����\;��
��z��)�N��o�=;˽J��>Dǈ�J�l���Ϋ9<^w�]���{)��O�ٴ^&�7�W&���C{�U%�ެ��W@��j;��Ⲛ8�H-/�:9o8���j~1�E���q^)�U�
lH��U.��VǬ|�Q��ۍ�^�dM���=�ᨅ���a�kI��D�󢙜���.&ސ��WgK*����т$�^�a�/�9�AXo�)�\0�|�Έ�A�G�4��Lhd��!�s�+���'d<ь�-/U�<i��5$̖~��&����jH����6ۤ�!�2��g}�RXj$�����b*�ѭx��@��x��tc���Ih�Ӑ����-ʝw���Q���\\�1�-�c�tV���rA�5���y�g
�x�Eo�b�=���阝�TT�ʸC~g��QW�"�E���"��0l�H�;A$E>^��֤�^p*{>I%�v�������(���c�B��]K��Tօ�b$���.�����ltìR�=)U�a���d"U��(]���/��/ߣȽh���9%mrq��D�M��9˾�>�;�GwM�9&�b����U�UyR3L�tm�b<���f�I^r�7�C潹�\fn⨠R���d
�Đt���~S�s%o��g�?��m)zZ}Y8��	���3n+���x�ަ����v�L�T��9/�r{�Fl�����O�d��P�@�;u����U�{��}>����y~<�:N�'[��]�I��X��^1����*�Sڪ�٫Oo"G�Ja��M��yc�qUD��Ι�RU�u��לּ
hvǘ���N�P���LY�U+Zt���.�f�9'O�u�*�ʕ"Qzb��PRĐ��\.��l'�7���U����)Z�XN6|�Nh��H�,K���� ^�A�i���y��~��s�:&�KD�v�gF������.�xknn�.rri�rw�6KQ_�XI��ϸ��S��a��J�R�W~l��-�\H�Ġf�K駡�P�_�eU��c'�KL��h��M���:I�C~��Y:�ӗ��5�M�B�Ѕ��-_��7d�fEW�F++���B=�
Nur��Y������x}�;�U�c� `����&��x��n��<U�pr_$�x�M���ϖf��!�ukr�{��es���

=�͢�7m�?B��H���ޛ1�fs^��n��j���h/L��,~��~�A� s����Du���:i��7朾��s�
�Qm��YD�hc���V�o��)�%q�ݾ٭��@ޔ�l�!S�YΎT%���p����4�Fܺ:��3�V�����S���*sd���Zu��e��}���5��c�l�)�Vi�_���R�zꅉ��n�1?�J脩�)�q �
h���Tې<)2��aʄ�t<�ˊR�:m�zRM�s[��z9�s��+�΋�Z�^R�yK�t����e�7��fl�3DԽU8iI�g�g��{S1�%�>��3�B A����?�Z�����
�/ʉ�"A:|���T�<���t�c��T��ÂJ�(b��Q�T{*�����>��Wɣ�B��rAe�Ʀq<+�/*����-/⃥���z���"�
=���q������nj}���c%�j
i�j���='�GeOY��^�`nzKL�k|��`��Xvm���H��s��S,W�+PQ$9�r�g��<V�@(̩lw� S��Sf7� >%���7�}�J�:	�m�}��8q-�;Fe�,�F7��먺m)�B�w�u����"�zps$�5h6$�i>֧-��˷�;�Jl�y��8��jxf����᪛�^�~���ӷ�1��v��!�����8]�Y�9$�r�ŴA���8�`�GZ6������zX(щB�!����I�R��˂����GQzƌ��8��h��?��J����2ѽ���|Da�%U�-a+��Q�4s�~�`Υp9�s�(�!����p�̦c���Vr�W�/Yb�7����)r��G�T�mk���w��gbB��$�������Yyo�:#H����l�-=�|�"ڻ�o�ۜ��0�H_����_?��r������k)��R$ݞW$^�8v�N �}�Y�|/
���^+F�!�#������n�4\o�Pb�� �(��rK��YO��F3�9,�AE�&/h"��wo5�(���^�QOeAM3~����&�d%]�y��[�o^y)��Z�C�pņ7vƹcbd "ʰ
���Aϳ�9d���������!bc7�AK���^[Ω�,�+^!!u)���W\��y^w��%+m��&Q�gnFCg�a�BW��L���L�$Ɏd>'wd��s��є��s
*Ǌ�*�5�vl��/�i
�/[5Q>�̃����*�/M�A����x ZB�i���g���K������A?���8���h�Ҩ�����.'��*�錳Ʌ7�/����� ��{}-&���uӆ!v�9Q��t"*<��]����GU#��&k��B�3^��7�ŎI�k�Ku����ҽ� �����!��?̠✇���]���"�;�}��G�S���󑷉��Nd�׮�>T�����ۋ�K����Q�E={[�w�n�,�"a��?У_�?��%��;[-�$e��y$�"8u����@W9�U��95Y�Ð�ψ�����Q�^ ��"V��F=�SE�����߾1�XcPo>Բt��z"��[+0���pCU �v�6���1�*�/H���r��嶝Y�1�g.��ԃ�*�*�v�R�z�U/WH�ԟMf6ڗ[�\��+pn_r)
�\t�`FrE/��I���6Atx����`NN�0��f�x���7\Ȉ`/���	n��h�@�v]���ɱ������N�o˒8HQrm��,U$cpU�kO?a�W���e�2Ǚ�o��45�|�e���3�F �0!֠E�.+k�w��R!ײ]I�b��漡RW��<Zc�LGG��]	Y���xIS����x�&U�H�ܽ�cD�����0��ĽY[|�ߏ�
�h��n{f�)<����OĆ�J`ʌ(Ec�¨������C������z�.ox�W<��w�Ȩ�$"�����MX�,�f�w�ν(����
5U)Ķf��������Mj�1 lxg�~ $�ڮ�u�<�=�Њ�������	()����Ec��pĄ[�JX}���t0n��lI��|ڵ��L�D��!ܵ	�5����8mL[�rL�1l\�6�ljZ�3!1���v:���åO�۳��Y��������U"��c{�yu�r����
��c�� 0����sw���C�F����S�i��7\��ߴ�ə/�+�Uɔ��������QԂ�|���:2�1�{K�>�a��y�N̈�!����� �)�0��ӄFR%��p)}�[z��Ty��X��n�ê_ma�l<�E��=�f��6��n &��A�cA8�@c4۩�,�\��2�� dq� 5VW4�����dU�y�b�B�鬋�M�����f�*���Z�y3�ʦ�t��0���
¸H��8vnj)�-��MB��u��)���]�9�9���Ud�d�F{�&��뿯��������3����g��ۢ�F��;#�a/DƜ�Q��S����i�1:��[�Mva޲�n���;�`�,��ckjG��D[�@a�`��1.�{�K��"w]�"8Y�y{o�$�~'�޺4L���I���`�HU!x��I�Z��'xg���T�O+�D[*߷Z�E�F�Z-�Ču.�r	���	�����{�	Q�e#������-����b���XN��!��������7_���I� ���Aǽ�E)j�0��*��c!�P�,�E������w-��DO�{k�ی":��m�LTdޒy���O����l�1L�}K��e�d ��AG��X;8u���@�0xeKPv�`���Pf17r|�H�:I�osw����Lr�����l�B�I*�w��{�f�6��R�P���ޘ���!��}ꥶׄ:�p.s^W�c�k�c5��9
�!:�è��A�)�G�d1#�v�� t� ;�bb+�q��y�������܊����Yf{�`}�L���G�L�ɜ�_I_��q|����0�=�Og����6_<'�p]�X9��*ʟ�$��v��Z xc�(�8Aߤ �����G�4�W)�:�?v���,Ԓ��8g+47�X����k�9��d�PTXOQ'��,���+���o��R�����xO.�Ɵ�j�]�l����G�_��ʨo
�#�2!���C���5 ���m�����F�ꁝ���zF``�O���B#V m���Y�A��=��(���$F�CF��Rb�`�H�����]^Z�?-��{HG]2�	�Ū����v�1g6�|7)��ǽ���>�s�gKAjn�>;Ӳ��1UҎ��.��|R>����@�Iۥ�~nR/Lf'5r�<g1@xo��5�����oS]��j�p���9�/�&�3�%ߎ�j��M�Z~{G��qUH;cH��\����X�� �!���=�͖�~���)���5-�]]�ˤ����"�����m�>Q�<4��Ӣ�mc]�/J	[�\j��q)���u��Q
ܐ;4����+�_݃��8����Һ���PU��T)1��R�P!�ʞ+��t I�_q�c�3lA��_�%iiQ�<F�>2/}�sy�zu�I&g�T������J�}�4�C]?8`�҆���{�w=O�Ç�� ej�Β��+��Cf�,���cs�a�����af\eN����_��Z�$���K��:f��5�d.l�yXwG�q��N�y��^괰=��0؜�]+K�����~FP�q`�6"�|A�{������������\|Àa"9���X+k/�1�L���C����y�ޫ��7v�X|~�F��1�����ת;h��zP���Ӟ�n��ZV:�n�+���&�O��jC���f���~�i�����.ռ��\�9�����a��.6i,Mn��e�G%S��s|��J������|,`8@�6p�B��L������w΁@˯X+-��+���Ag:<��p�1��˦��Iz,��b��U������'�}#�R*�O�P�\k�i8�P�2�)@�����9�_G�x�ѝ6��6�����2$n�N���[��ē��X�Ya6#6	r���qR'"0W�9�r�9�]���k�Md��j*���"��]��� ���P0ȿ|��jBDjC��;W����!"��`=Kp�pC\I1M��*��^�~�KD�zI��i�7�6vAO`�E��Ż��,C8���|�C�A��R�2��.�� D��W/�25���e^s��0*�#�\��e-|쓹w�Qb�D�O�� �T��22��j��>�JioA1��k��n��׿5�'NT�/ic:\���0�a��ߪ��b�oA�Y<�$8��!�J��o�̪�M54�\�5�F�Sy��t���-"��jH)W+
I��qS�}=[�L<� �Ux������B~��M���}]�|�'?��y���V�E�3Iךub,�8o�W	D����	��T��z'w�E2�aK��!߫b	��I�v�=;ѣn�tr���dtgS��yR �Ȯ�j��Ne=[�;h����z��>��5�����Qy���\��c�#�P�z@ؤ
0���Z�'�bf�X�
'vx��lY`�:;���8�)�]r"0�Ō�溥w��b�{����CG�����y�o��C�e��l�H�U����R��`����N�f
\��ZT�"��.��!MRh��Cs���Ə%���"�y��6�N�χ��|)�����o��U�q�U����'��;�VGn�]�C�u���f�1��_�K{n�[w3���U��
-e��oAoĳ[��Q}���5XF�S�/����J��$����9����s��$\Z���8��㏆�����#�T!#6��g���K��N͔����^d�W�h�U�;���$Hc<h;��#�ESÓ�]�#�rP�6��lM��|����[qg�8��NoO%��o��j��ՠ�U$P@l�q1�4"~m@㏣�I����GL޹� ��ϭ��HHE�98���?<}x�Tu���\��P�Oµ���\/�hV��;c�l��<���\����!��9��c�<d:~JFi���aL���'�U�W/��&QD�<��į1
2�`��<$�XI���������z�vp����}܆�5[b����R��86�h6���6M��:(��T�A�~�R��?Z1[����d�GY)
�R��S-���'�s�s�^C�p�� �����:���'��S���7��{hM�,�q�JNe��?zB�с�P[�%X>��z��
T�P�D�^��բӦ
B'��2C��g��ČМ�l���X%�>ۓ��zX����x&&F��������\��2���S��yV��*n�DV��
�,@�r�Y5�ټL@D:��������P.�6
��Irl�8N�
v�\�����
�#.�˭;����F��j�t'���1)��9���A{.����]�����i-hV�����Z@�25b�|,�.0���4>� c"_vt���4�����YҘ������kT�&ud �YI���H�����J$��N�N�g�&3�N=��uBh��! ��_y�E�w"�C��(�.g��/�xM\c���.���	����t۾������r��sV��s�N�Gf������z��֯�|���m�`j�#MJW�J���1Ҽ 9�����̑�α�SOy����(�.nŶ Ϭ@�xd����&����ȡ�U#����F��c=�E6��}��D��h*��P/�䧄2M���Dj@
����s�o=�1%�Y:h^o��7EX1��^q�<��)k=�Ƞ�K�Xz�	%R��𰡊T�X�Q6R-�/��3�A�	�A|���2����!�ώ�����3s���#����6FZ�F5��1e]sJF���r2�\rh��r!�H��N�'��!�vd��׷��������1c�|,co|�Թ/��C���4���¯���%�+DK�0,��4����e>{,?���W��&�"�D��3�G6�����d#k��	��0��ܫ�n�O�Z
���2T�K,�i`����贽kG`�Y�H�Gs�	aBbF��V*M��s-e�>Z�@n�,�fru�4^�bz�?�C׍�"�:i {*�(TN�� 0m�Q>9�'߃�^�bv���#�4>��՜-Ȗ<32u����U:��^�"��/��W��K���F��%~
EXN��q_��B��g3�g.�89���mc+�U�<gi�MwU�ld�g��a�����!{��d����p�58�mfA�����	�sv8:�EW#���-���h�.�޽�)�ճ6���u
}��Վ̿\j�<����m���a��(���^hZXI�v��Q�^�BY�mo��x걣̤a�8� PH0�M�
����z�g�)����;�M�Ȉ�$�Υoj�ï��Vѳ*:oG�n�L2����:�!����Q/>�]�1Q����bes�t�(���-{��i���Np�p�O�On��v�*�{.�K�h����0�6�jh�t�(���{�zu��]�t���׬н�v9(oW�M*�FU�H{�^{�ݖ
&P������1CSy�J�UG�̈�q[�.֠�ةWN0�3�%���D�nم�cr:�2ו��M{X���T��T��O"2��@�Dw���C�QL��%ˉ�Q�\X�\K:�-#+�OwR�I1���Z��X���.�䢕�t�Ԋ"��EqG���u����P�,4�s�G@�;�p�UL+!]?�;ޙ[%֘���e1��ߗ��,��@�V4�B
r{l�����<*jz���ȩ��O��-�12����9k�X�)���fױ������O��\�'�� ��t@M�n�G��	M��o�+�t��g����=!���#�R�[nM;A��~�Y0���I*i�K�er�{萞�Q�������(B��hO[��R��{^��Fʦ�X+�����h{Rw-mm�'_I����U���c<A۔o]� v5�}g,�ryS�qS��k�_̅��L�����v+��H� ���W�,�Z惢{W�H�������X�J���X����j����f�Ic��?R���E�@�l���q�"8�����8�S�����K��v����a�0(�8��	g0�xvR�Ł�Qϛ�o���Cbr�ʎIP�b�j+�=	&<��#c��_X��B9��<������} �S���K��_N��ר��v>��o���A�a����d�t�0\O=Uf�%:G�k�N�52��k��n�s\�*�Z%-��4�.��	_�:�Z�Kӎ�v(��T0ܳd�N�WStƆ�$�)�!''W�槽�V֑)�e �X�����ɲ��e��x����F�FvMZ�y�g���IZ��/B�IB�R�]PEj>�j|IRN�exO��DZ+>�f�L�V��X���=�T�|��?����� ��Eo���]Q��@'7��i�
��j�?l�q�����?�w��"�� C���<ԯ�XDϫ� ��|B'��@ˤ%:�]#{sԱ��jV�3��ك�&��	r��������HQ�V|1հ��^�T���NN5	[��e[���d@C��MI׻��&{���i�!E��C����:��.��8)6w�[݆���s�v����C6�(���bZBjN,؈�'�Hub�\r�����=	��6�z��5�غM\zXU�'�3Cbk����7?ve� ��^�:����t)�a��
Iҽ�=$1�bj���|+/�Sh0�{��͹����qjAS/���a|������E��>y��%���}͂�kf<R�"�26�ߛjV�
<{8h�R�I���,p��&�~�O('��$��!M'�-E�zu&g�Aľ��e���Z�����(ąO�o*���
h���hMr�z���HNn�@�-��`�H;�v�NwIV2�꜂Κ�q��K����%���:�!��C��q�<�`�|�~j��j�&!�&* �e�ꊾ����BԕD:�L0�K����O\�=mA��b-rGn�L1p�@Ir�� }Cé��V������#����t.	 ���wb��R�w����Fs)�ؘ�S�r*<�r0c��d����ug22er���bL�m�r�[�"�N��v���>k ��;�u�N����Ki@e�����Ed��W������x�s�Ɗ��4�����D�5Dߔ�[���5!���j�ab���C,����x�+NK�xI�;D��mVv?����1m�X�Zp��/u�0�)���sd+1Ze%)[��������UV��F��iU�XƋ�T]���r �	p����e�ޓqe�A��q~[�VH �ͭ =e3�ޥ�9��Sz5�!`r�'v� D<�)!�+��*.#3*�e����8k��dP���N!�s2:@�����k�������.ͣ�|χ�����C�J�E�*��de��O��|:�+*�)%�i�����Ӑ��P!T�gWn��}�y0�P�К�����EC��M_�!�$�}�!91T&�yqFmL9YX侮f�5B+���<�F*=ߘ�m�O��k�sR�U�6�����´�h� ̓��ط�f6�˹��0^������{Σ�.e;G^��<������|ԔWXU(m�S�Cv��I�3YsH�!��X �_�4bhXR��f ��SON������_;�s��m}���H��m�4��2��j�#�,]�պ�EB���Ĭ'�}a�1I����9;��c*��n�=$&& ;��}3�k����q����p=^[��[�=��t��wą�Z&\��jU��� ѺL90C����j�M;����"��t}-�ڔ�D��Z���� :���]�:��d�gE��!����ba�51�j\u�4�K�Ŗ��<r�e}�_9A���{\iM1~��٪m�"�&��>���f�u�=��i�MxBG�m'{��Ts��u��B�껎�5�I)��	AY�����T�gJ=�i���u�ˎ?KR�
��ߌ�0��zP�)�P1�@���s��Q��P�E߼��jN��5lA�Zu
*I��hTpu�v�[k!�7��H�eD�~��-]y���'��:�jHfE{C�i�߹��+x���`PM#��:�2�tG�N�s�_*F���
qV&�q0�O��V�$5U��`�#ğ�Wp������A�Ί3�����4������t�p���Z� >����-��9魆¯���m�|�����~��&�?f�?����^�\��g��A0 �O �����d�җ��NC
�d�b`z�4���1Qt�E�Q�j��HT�=���]#�$�C�+�O��PΩ�� ck�rSX��BJ�/X�`V�B�	��.�	1�����n=DJo*m`v��}�b���n����ZhuEh~��zg+q��p��c�6�ۏ+|���ׄ�aj�vH��'�
��DBO�ڒg`����4L:���>����@�_Hu�u��̳U�Q�L~�d�)�c���~�2%�r0DOw�\�qb���Uw��C6m�!S���z;���ƀ��4d� +�-��ޘ��	���2���5��2�O�����Kk���m��c᪗4�N4��W+��n\���Y�g	��џ|?� �OuXc���_�L2"u�P�[�l��=k�m��59�:���}	/�D@� ���-i��4���4)���\�u�UZ\A?��X����������Ux�<����J�+�A�*��(���8M�}r���"�v;�CQ��+{2��
򇁸�]<1�iGw�?����h��E�"C��%�݁j���z0�".a�*0\8�,|P�Ȁ���=c��N�:�.��PA^��������ʍ����#���hP��w�u�N��9)������N�G\Tf�x�g�Ñov�m����E���צ�=���$��HC�� av�1���I�`����*���E8�K m�Sb��n���!�fB�S�b鞥�xe��w�c�ebª���}�����Řc`>��<��(�9�㱵�l� 	� ��{�>D%��sV���sN�ր�h��n#�e�[h�U�QqV�z���C�.�T���e���/�¯��AC��Q��Јc��(a:M�e���R��ڴDb���pĎ�v���Tw��W0|���)ud���	*O��3�*H��DetKS��ѨG��t=�2z�"O�r	ykF�T�(�x
e�ݶ	���ݬ5��0�,�`햅��8�2`���S�NQ?�9p4��cu�^$�z���Ut�����Z���@�;���'/�<����h��ɃFo�3�������5����IQ;�� e�]g�s�2�\� 8O^���gc�o��s�<�Үr�dƸ��dpFPgb�"�ˆ\D�(L�9c=�r ��������	�B�S������B)\�&3�^`}U~�THZ�5��o[/�9B<�����Հϑ�:�7���Wȥ=Z2On�V�����J+d�5�%'� U����u0�p�`���yS 6���ٵ9���B�g̚�
�o��2�(����^��DTo�~�kF('�s=��!y�������3\v��f^����y��9��C6����I������I�!$�#Р�뉌��x�%pC�G�_Z��}��;�1t4/ks/2#��2ah��t�U<�dӟP�F�|����XQ�
����U��x��x6_��C�`�J�
��%z%��5 m�a�t7��;�wl՘��p�sft�=,�6�4�H��B�o�v��S���B~kQ�| �0�1�@o�%C��O�R�G�;�*�v*r��U~s���]I���{%x-x�拓Y&�_�(�B�/4���.p9�H�H#lU�,��(�~1�8�LwM�>��D
�Ҹ R+.�,[�h��2����S�J�:�6�I�5v�;�2T��L3�x�Z��?��ݧt�VXv��<��]%���!��qxl�UT4���y��N�I� �[.������"	���jK/-�y/�."��Tu,��x�f����Y��z� �g��˵Yґ��>j1Jp��a}��(�UW2c��<�o����I��XMHM"7޵��%}��%�.����KF�I�Ԛ��d],��ܼ�K����H�>-�encw�7L���@�r����ư�_Cs�{��yi��X�r��I�J�!��*~���y���*��y��zޝ�OW���א�b�����}k���q��Nб�s�HB�Fq�܇B;�7�'�h�=� ����f.dBJ��ϴT�	�q3Dwo*�u���X[9���2�ZM�΃��̂���F`B�9
jX����^m]Z�I���6M�@In��X�"��v\;%��YK M�� E���&�5�5b�l���m�ԃe?_!�'��,'��<�3u���Z��ծR]Fz�`uM��$K���7MOJ��m��:�T��2�>�a?�4�_�o���?b�(����p���1ެ�\�L���M5i��x��>������h��8��qG��KυHWO�k65X&Os��s�ׇ��j�Ү�����a(��٫
Q��y� 6og&)�~��N���`�ϧs)���`O��4�7ֺ��ye;�<��5���Wߖ&�ɷN\B�S�$���Mv���3��tǝ�cԠ��z�>h�<���^.�r��V�̤i���_�'}��P車^�Lh{x�޻�	���u!���`�Ҧ��lH}�!ҨJw�'T����8�ݴ�ݮ�`)$�/�"�@{���z˜���
y/�tU`�n�v;H��?`A$���|1�D�aQ#Q���3�9�F?8���?���5b -���P�%p�Ta����� �{H��be�z{l�p���e�'�	���2�H�L�z�+0��b��$y��5�yب։����"��r�~bǖKO��"�z ����s�,�⸾�F�3,��ڕ�(㼬��4nC��ϫU׊@+�_w��
�dz�� (�h:����-�s)E6�Z�N$�ū�������"�^x��/7�4
�P���z@n��� ���z|e�fX���;�;�~8[L��;�����Ur&�o�������j��C�<+2@ڟM� ��\�OD��Z2|��^�P����m <�f��vp��_����s���A�_���ˢ�����\�C-�\Oݓ�nM�����}���)3p_��p�h{��:8�[���*��r������bh�%F	n��w�]S�3O��h���ZRǗ�`�A ��=~�z��%�k㞉��&��AM��@�����\�|yєOC�ѹ&�Dj�r`�h >zZz����<���H� �c�{�nn��VH!@�0��Z�`�
�rV���e0�h�[��0ܯLϻК"�sf�i��c���#�;K�8o)�-D��V̶��O�z��U�z��Z �k��3��8y�w	ͫ�W�e�����+t�вU�h�X��y�Txb�bA^P��81V�S�_1����_L�e��g�`I���Ȁ_��asȝN.�	J_g�L*	�,�v�f����N���V�>z�s��x���cr,�W��S�zz��4�#j`�����l�&��4(��}\�
�S�=ٞE�u�m-jܸ�����[�%�Ѓ�D��0�� �ƭ���C�����%f�M��*R�;w�N�ҁ� �3���p�b�kl�_^��<��ń7䵱�� )��\��[�)�0�B�o�&-76=�OԦ0
iT�6'pŜ`���7�����@�Xڟ>M'�}H�b�RXj������$��i���䒱�Q(��n�Kt���ڂi[�٫��ث���T}X;O UU���>���{R�;B�̼�F�B'c﷉�s��#���0���2�=��4�9�\_�6bEnj0lZ�4�xBZC�"�X�`V���s�U �F9�>������Ȗ�v)�a��r"b���+���n�:@�Ic��mV=�11z)
o.������"<_��~d1�]z	����v0m
'L+��d�1?�~�Yk���~OԠ�x^+~P&��Lo4}�M0Ta\K��k�3���k���g��e�/�X4*ٲ�0��=�T������|�`є����|L�	b��h\ b+������)טV�Ыs�C^]O����w�� �	y�.�;@�pt�U)ӳ(6�a�1�!����R��pn�z�U ��+��]�'�w%|�9�����%�?�:Y��,����Þ ����3�Mx�d�]�.e����o�df��_���x?5��v	};����0^E'E��)<V�OA3<j3G����$[LPI��`�~��Nrϻ��84g��s|[�l{ �pʉ��G�c껐�ߊ�t+�XX)��vqu6���h��r���sc�����D�3H��|�C���i	�Z��1���%�I�싼�K�}��~*&@~�F�qf�6��:Xۼ��I�0|�am�zh��=]������7�u�.�|�=��#��=�|Q�g!
����M��b�|�Z��6kAC��Qg��u�M�^ߌ8E����8���rM���9J"a$[�qI"Eo1�ڬ�^�#6�?�  �ќ���kv�9!݇�@h0��*��#�<����Fb��oQX��0��Jq4˕�X\��u7�Z����X�KK���B���) ǎ�t�I�X���X��<���ae�F	��~*8w8�dgg�UW�蛩D��:����-�Bhx�܋����"~����|��nL �}n(�D�m�ڋ��#��E�E1�W�p�|��E'J��e�(U�6]��O�yY?r�)HZM&�`�J�;#�lV���45)If]�6��q)��kE-ꘊ�o���d�&�S˜�[$��?��^�A��s��`F��1���v����N+m%�1f�@a!+�:�k�Q3=�o�s�]��跞r��� H�����U#CP��u��|B׻�pл��iJ�>VT{~�=�Yx�K[B^�����6��
�Zp��#/���/�	�5�-��Qs�ъ�o}�wWm�T��������c�`�1[傕\�6��eݫ�~՘����؉��n��$(�/����a�9)��V��ԭW�����a
������똲Ya�t��8v�;����f�r�ՎT">H���	�K��.v*D'���G����/�A�9��h����v Sz+��!&��0q8܁�6���,N�g�e�����Tڰ4��[_`�+�ȚGQ�}b�b|�4e��[��V��XB̔	����]C�Κ	8��K��C�>�$P^���;�!�����o�M�/��aU�o@æZ Ob�?�$f���\O�i8�*"�2��bdt#�<TQ�C�(:Re3�H�#Z�HVA�~uq�~5��Zwٌ���	���L+d��BЦ�b�{�Z�����(T��gN"��)O����/��y��_.���N˅�ΙU���S��yb�M?{�tN�4��!!T�\-��{D��ӯm���XR����X���s�k��r��sY�%e^*9��4�7�ŐE�֡m=ڞ�`����h	&�U�[�Kv9Ծ(��7��xp����p����C"��.^�kI:�'�'�͛��Hl�Q˔~Lz	�y��3�� +]�yQ���`�5���#��gN���3Ƶ�h��j��b����Ň�t&��>b�5�L�ql�������	��\"ҳT��H�>Kq�m@�v�!.y_ru�MS#P鿎Ç���[�G��WPR8.Cģ��%y8ٌ��a�/O?���l�g�@"Y���ؼG�����RF�����j7��ލ�leH��B�&�C�m)�1��P|�����XM��?�˨˼��_)m�s��c���6���3�Cx>#g���|�6ы�D6���q�~!|��g'(�v20�a�t���bo��tBS���Vt�_�Ҋ�.AR�{-I��°ĳj��>�	1P�r���_�<���ø���Le��R�WUs�޵��~���Ǿ��b�&��v,�d�8;�|W�:S�-����/�	�H����m�:a�FDrAI���'��'���A�h+^Y4��?zq�A1X\2��|a~�VP�o�A� ��(�}�ܧ|G:a�'ee��|��J<�3ab&�W��2˲h_�,)W4�����Cuxپ���	�*ST.����~�ɏ�idJj>K��/ˏ�^�i�7��h>��S�O ����`Ӈ�G��ٲ����z��3>�\�RxP���Շ��`�Y�|����N�1^�M�@*������Cxc]<Q����I��(PW�"^�)^�g�&���,��rȇK%�Β��kZɼ����k��Do�l����ހ�#�/t+{H,*g!��_7a�r��o�O��?�Qʙ|D!H�}z�T�P��3����X��������x���;jB�W5�e� �tO�=�n�_@HN����2
�B,��SB���򆮝�)	��U�ٓi�-�x��Q,��.3�+cs��Lc���0>Y����3�x;���{<J�X�59s&I�;�#�g���1�)�ִ�*�^k��Q��m��ȳ3��M��#Mđ�"���([�"����1*o1�~>r?����n���j�.���٠uz/��\˟rS��'���� �h�	f4p�!���k���ng��/vT��a6�^�h,��uE<��<�9��I9}������*F�u�ƫ��rt�p�2	8��K���9��Pp����s@3�b�>n#=��F���f(4B�,�M��c��$1 �çiv��u���Pc-JG�u�\.��oI!�(�Ұs�G�t�z2��.$��7����	1�h����A��F�ۥ<<��Ԗ,)�pO�$z���B]Y�Y�ٱ�C�#���A��8p�|�G�J��W{�u�צk��`�	>(!I^Q��
aRz��0��@c�b7����4��|���������7?�������m��`�v�<7���^���3�lU�o�}rw��i���� ���M��-����Qޤ�|k�[�����Z�X~U�K���J�O�&�8���_���F�.c�n(��'ߤ����m�&����{70'��e/�"�㦭��T�&~Ҡ��l�Q���g>�#}�����S�`�K,�I�����4����XP[QuZ�vN	����ޱ����)Y%4�&��%Pޒ�C ʩTՈ���%r���|�s�ZZj�^K!8E�
�;;+q�9�,��C��9d��60:l)��v��ҹ�..��8�G�?H`n�$8V���yY���(���+��	^��"�	�ϧ%�����kH�����߻��]Z�v����҉(xd��^��[mo��*m�Z�����&A��]�T�E�%�S8P����MEffCʜ]�ތS����W�3�5�ġ� 祮w��`3;�������jf��@K�<�K���#{ƃ�z��&����⭜����{�k>,A���lAq�{?�vG�}����A\�A�O����3C�i�jy������4�kUո����4�^��x���L���m�f���O�ӻ���7Y�Fx�"rJ��v��ϥ�WbIK����~L��)���rq���,srB��ڙO0�G�D������U?s�U�>$�d8�\LO�����o�՜{C
���oyR+.�r]`�*&Pm2ي��9�.#G_'n��e#uvb��_�2ބ���Z \ ��pB�9�u�La/�R�m������(�	��@�f�K��#������Es�Pt+������G��e|W�Z=��ܸ�k|L���3�@�� �;��M���/#a��=S�p���]V��9��>�U�!��H��o�.)s���)�I����A����~�ez����~�+L`8>U��?MD����|S��)�-X�^pѦ����p���Yp�E�1G12XX�QP݆W���e �������gT9h)��K=J�r:� �e�r�}������������8�d���R\�҆����+e�fnm�E��o�~�F�2�r���IC�ɛv-mqc{��	���&��/�#�*۹�J��b=Y.�|���$i	��}[��0��I�F��]&�����B3E�����m��N��ϴZ���*ղګ�&���0���O�m58��z�y�_S��m(.��xYy��"*d���Iy�J5�`��T��<&W�k-���%*�[�*$^��� �SU��r9ɱ5�g
,���7<A������N���O�����c�)���u�,0G�|K�D0���q�a	E��y/}���}�E��	��L��� k�P��I����E�^��#�7�}�D����Iie`G�͚� =��/�k��({ `����仕�ʙ�i��>�$��5�ol	�e<���9}r���,�=��0fEV�op��lC"Lβ<q_�k��\5R����ޡ2�U��!��#g�x��@�7*�C�0���o?�r�6�$��j�[_�'n�a�IN`v�Kg�,'�q|�`��x�Q��s2�in��dL�a��5�"� 	�ߚ��u3z7��M�cZb��:~�e���{��v���(�%��
!�P�qǮ���d�H"�=�Т�Ν�FW��R�pd��bG�P!|�9��ȫ�傸$�d��}�O���0��;�'dS}���(�j�\�P>EPړ�G�/ix���7[eE^��������B{�n���Oy����0|{ۤ�y��C�"�K|��a/�I�̐�������D5ެ�܅���eN�T�eH���AZ.��.��M�%٭�q����J��*R2����3�Oa���Rd�քM.7^���;~���m��d�*_N�Eb��2]��\���K�Kt0�M͒���;�Wѥ ��~�\g��$Q�"��'֖�ፐx� �LJ��?��N}����W)�YstDl�h��8@V��]W7�5�Ѱ��8�28D�ԇ�1�v�cDb���.��0��p��P�9���s?�>pڠ� y�j��Q�l��kw����F&���!�-��y!Tܚd��\���nE���+��Zj�x�/�>Rv��=?�Mg���<nҪ�ju/�B��Y��оkcG(##����Q���3J��#X|,耿Ɯ�:��wlU�K�(W�p�"9�j�V7�H(v�3HW~����``�x~l(���#`�V ���i�)�)M�` �ո$�.��>g%��%�L!�x��+\����(�q%�>X̤����a��Cl�*`-�̗�z��هG���p�>�-��I%y��d��>Y������Q֢�⌯i��ǈ�;��R����y.���4/�y�5<w}�k�&���O�\��*g����� ��*M/�sL~#�A%6�?���ׄ�D`�T"�싎�r��6a��cb1e�$�|v�� � |Ig�o�q]R�EN�����j4���p0�DN̠y�J���fd��\�o�E?n`P��B�����< y7�2#�J� �Hw�j�2;����͆�Í,�|U�2x0�R�+��L���n�[���)�\x>�q��0��`�*	��NC��폜d.Q�o��l�GqL�v���X��K�TbZV0��!��g<Y�dT�	^�2��ʧ��y1��04��\�ڊ�H�0��T=y��@����:�ɹ�9q��6�A9^'{q(7�(���WR�=X�	���R6�|�C�����`��C�����d ��A2,itj�;��W�Τ��)���u�cbɄ�H6��gI�|��>��6����W�cGb�؅3:������(�"V� ��5�4�yl�������3	�^����Xl���T">�_�~�}�������j��o'�x~����CE�a���tF���6�w{�R��9����9p�j�̊���]"��@�Q_��hړ��LF�@��P{�6/';N�����r;�v��=���+���q?�#kμ���),Q�W�fu��PB���=m)������g�K	�˞�	�uD�1��l�����PG��J��g������^�IkAv����թj���অ�?k�_�՝j�Kue��^0�_����G&Cs���	�%U�s`�Րm�;E��gܯ��1Y�� �Ok@�ã�\դ���XC�mn�ƳM˵�'V6�]ס��`��EIq����'A�	QL@��3��N�#�u�?d���XƎӹ!�oh�~+�p�1/�.ͫ|u�51��z&)�X�� �m���K���f6M�"�jtEm��}�>b�������{������g[8�'QA��HeƊ ��6-��3�G����a�DѲp�od���XZ��e��&�I���&b��E���q�}$h�9�}9A1��*(1v�)��r�8]ş��۴�տ� F�VJ����w�2��f:�	a|0�j��	�FD��|��K�a:-)�y�.�,c�s�Z�<S��'�Ь�� ư�+��e��(~[4>��/�"��E=n~��Gs -G%��b�.,�S�)\��.Q���"���J?ִ�ѧɹ
���|-�>7�[�pu�G~�&��(���{����r�xC���~�\�9�IFR��ČP2+����o ���ra5����*�z!��~o@[�˾���%/w��/����ӡ��;��'�t��H���R+v.e�x'#B]�����*��D:�p��Ӝ$�s[6wAl�ڀS���!�6WSe��ր/���W��͐��#��^i��~Ӻ���p�i�Ө�႐�h��8�壼�ݲ����,�ثk�1!��[Z��B���(��@�e/��r��#�^ٿ3��.x&l
�P	�{O�'��I�TH_�]G�J�F��O��߰_hC	M"9]fI|>��V�"�r~�b��n]B�Ef���hr�P�-����Q�)�|v�xFY��G/yJ�x��$�c	G)N���[������eW�`I���� �mZxI����z�E(`b��Y��MO
Q<c�����"�a�9���۾i"#���:�@��~�y��v\�vx�GwА�<L
j�V8��4q�d�I1�X�HG��ԯY��f�A�\�)��Ӓ�l��]�Yȇ�;zý�+}�K���`JQ>�I�����۰����+�˧�׵PBM�wR9�k��1��^Y�n��0���$I�Qh1A6"��頩\��m��Z���qFY5i㙑�$./j�0�n[�]�o�`�B��JU�5��	_y�y7O��@�ھ�|B�����}����x��y�ͮ\�i驤Ƣ����� �jz�͟�h�a>���@�-K��	W���RP�5m"0���ʀ,~� �@c��NP���4�S��+�\E�q��BCp�~�'�$`�H�_�7��]��}���B����h���F��g�&&(�d���o㔥�@ǴQ�N�����R���uP�B���������Yt�����&[�h����j`������@,e#p�s��ͮ0*����^�5���oq _[1���A�<���#V:�������*�?�y���w��n^i�|�<~�E������C�{8������k]��2�Z*�3w_��d=�q��H�O'�Bg�!��tU�,?���1=F.AWUc�`R����4c̀5W�J{������:w�z��T�W���l:z�m�7V��E����I���f�pVD�.:&��a�6vb�+�Enڊ����l@+���S��xi�����"LeѶa�Z�A�;?x�;0G�@��w눉s��5�~ ��([�>Ԁҧ�P�|T��pJ6��^pX�o��45ڲY���T�Vy�wY��{�O��`�{�h�!Q�������ߒ���K�@BM�x/ۍ������v��l�Қ�����`K���H:Y �S��_)�Dcd�vi�kY'�����94gM!��13���Tn�[u>�Y~����
�}����H���Hwd��7�r@ۗ�O��dO5 �����+��J@��I͕Cr�U�V�0\�q ����B���@��+}pM��%`|��oL�<��D�Es/M�%�U>���Np5ӎ|>��¡d�����A"��p��0��2��	����R�<�bl�yD\���D�n�&��j��g�<0T���xY�Aqg�Kޜ�mb1�ݱ��% �'��䐜��d��\�W"�3�%?�$���)�T� ��}�PR�m�"H1�i�aB
P�7/%�q7�e��]��ӆ�����L�p�����_V�
�`hEg�R]�j[Bi�;�����l�(�x����8{�5��e&�]������H�r,�
Gi��V7ko�xc�{7M����-$MF:#��� g
gTsW�C3J޲q ���~
�����X�&���I�WE�k��YQ䑐��&=�Tq1� ȋR���R���9`�.m�;�;Yk������)�!c�?��+b��w?0N�ʦ ��J�����Y��h��۠U��C�Z9����E�`r�.yH�`nS�u_��䴻,oN�hY-9H�~V ~�FG���1}!�lA Q���7�(1[)��9�@ �/�V�y#0:K���l�P8j
o��mcr��ڷ�ah�^�V�����:�C�/�3�5����6�f��QH�������Vs�l�!皌%X��|�ִ?��ϊ�
�� �U9S�r����#іq�C��{��Ǿ�*�ths)!g�mI��~v�W4��\S���K�~�<���"�%1�4�T��k���1Tv"Q��9g�^�}�߈%�����R\���c�9�hV=��ˬ��3�����&Iz�:A�00Ǎ�9�M�F�&��P�1�&.��۲��׵�kQ�ƻ椷~��[g�����y�������\_�3֧תQS����N�1�\+e6f�:��:��3;님�>+���ah\�;��5R��Kܱ��Hg��>?�0�H4B��1���Cg0O�j�+��zN�����"�
>��e�d'�r�(gu��Wdy/�\N!s�n�XwKTY7���
�՟ϻJC1[�[�>�UR'��ۉ�%�z����m�]{��G}�N��#G��2b��-��&����89���\yŧ$�̴��0�ir%'Č��Ψ<y���^�HF��:4�N��xdx9� 8=��p���k%&Ǹ-Uv���}-٧?A���ܴ��������z��g67����1'Tw�{�<)�qT�.1���-�BUy�e� �W�<m�ܛ�Y��
.4�t�Xso��0��ڔ6Y!�W?y�����Z��{[�sێ��ʃrq��{��z�1G�ۇTV�4 ���H����4���P>B) ��.��m�rK�TX��a��YޥH�i^{�o��(� ��k�J՜��@��N��Z�H�e�R�f��r��.�+��2�p
��L�����"Q����*N6>�M��b�-�=ټErH�1��m��%���V���?fI����n{�E�G)g�(����W����~�R���dh�K.����Y)�������K_lU�")�2�I�y<�p,[o��7�}�7.�Lg�����Z͐0�ҭtZ�;1Mn�����^���dy�-�����;��Y�9q)���f[b���W�H_H�^���������	��x�Z� 5H��#��K4NC�s�c�M<�>7��S��r=]ΒW�D��	�E�����HbZ�%M��a�X�����|N��6K"s�����w7���l�a_�a:��9x���]Ŵ5ծ��0O��m	�}xX��$T}b��x�@�7ݸ{f>��s�t����QRq������j��m��>u(���"n�$��2���P޳�#8R���0BI$�[�t����W����P���7m�I�NHzz���^�EN�_+v�z���7�����E�]j!�,���S}So��=�L$�A�I�>a@�	�&���6�_9�UP�E|�2,�ZsbC�9����(�����l1���h®�3�W_�Taѷbz�����v��fo�@�`I!d,�x�duc�2Y���,�{I(�P!��X0����V2X�'�ʬ��xT�	)��〜��x2����k�Vn#��I��M��G�5b��-�[���C���TE�2��]�!�>��Pʯ�'Zn���I�&|���U��,�γ�� 	�o%�;�>_��5 �b+���� U ��Z���t��pB��4H�<ԥ��N-@�I�x���ؿ3��s�N��gT!��[���T�g�i��e=L���*?�;�1`@�$��L�4@z�j�|�ތ�	&�s�ܮ�n�TL}��7`�L[?��m
�)�����.~w�-w4)�$0,�����4"���缇�e���rh�ΰ\�m3C�ȿI��ۣ�VcU'2�PHӷ�k��s}<z�H����{z��kP��?���R���"���ۀ�!^9{��h������_̌_q�%h0ɍ��� (��9�0�읥��jC�N\�PM�ڃ�BdŎ��G�։]��� �����"wW��f��v��svZ��Ph��Bq;�N)��&4�N�<�s��.Y�MYGX��Rx�nZ{,�������|�ɝč��Jr��O�|�J,!Ń�g�+	��o�HiNQ2�fP��ˎ�1�MD}q 'T�,�.�k����XcX����N,��A���6�aQ�誣�H�j(#u�-�y�0��4�E0�H{=R_�&�ߎlm��A���D��V�N� 2��SL�e��O��(�/�R�������g��.�����?��Y�_����fc� ��c���^p>+x�.G5BQ�Y� ��@7��r�;?�J�DZ�|\Gl7-�2|V̽(�1��
�C~	��0h�f�bCxKZ�Kk��рy��E�8d�0�;�V���G�����|٭�aݚ�T��n�N^�
�+�X�~!@a3<_0㠹S$Cy���ݹ�c)�T�K����Fc���8�^�L�`��.�@R���e͍Z�,R���.l%bR���)���h�>r�S��,��j	�6�VɍY�.Y��}ځ�^Z��<9��^��`�827D��~š�6	�Ĉ�I���ٞ�g<�v)�Q�iE�%���7��8���)62T������|sq+�¨x>򙺷�a���fΐg)��;Vt�yaR��A�\�Jrr�K���k�R~�,JR`M��h0p+�o����u�)�r�XŁ����o�Ea �������
%�;�ώ\5�|�*3����_*s$��?+6���d:���y�ߑx(�X�TaD2�e/S�W��JH^0P7�|��^�5o�Zk4��l6c{��8y0�U@�N��	�#�"�{�@݄�,�S�0��}���+80��P��Eɭ��`�
!-(��-T�;ɼ'�A��4N��*
i��X�ce�B�o���[		�4M����NiD5ƴ��\��yH專c�j�Uł���o��7��\V@&�{e;���(���'�p
[�v%
�e�.T���E�5�Pz5��,��vu���A�nY�,��*-h48��
-� ��ko����g[�~�D��m��Z��<5�@M�e}K�&���cgKTr���oc����x
&K����_qՆD�{���$�ė�`��)�@�(I!u��i�/�a1�����~�-���4M$�_��.z��HB7��-͉#q���|Omi\=�)D*_�:|�H�1h� �I=c��oI=���ކ�����^�tz{�Lu\@o�Om��|g}�-o;�B�@�z�P39�<$ɟ�{��Vd��@�`i��̕3�9y�C�x�@�PB��ݱZ�1u��}HT�J*��?Y�隇��V������5�i�["��DX�� �E�U��ɍ�I�M(s:���&�q�=^�A�po��4�0��3�D�ғ� 1QB�7�W�ٶ�|_	�-!�d=-S/.�D���� +�ml�H'	�lyw=���)����[�N���lB���� ��G͎�Gi�'I����!��Q����*�ZJ��^~��U����"G5>�q�,�����y����$Ux��Y0�=
>B��C��S�Q�p9�����C%��&;�}Cb�Ϧa���]L��;�b�_�Օ?�#�:�bܓ�
K[L�O�S�:��鈾g _sM��;m'Y���R��;�:��*�S��B�Sy�y!ѧ�HY�hl���"�1��u�_;j�-p(�=�����ni��,<jŎ{��P�N�`֗K����(3�G)�'9Xi��v~��x�B�� �>3Ǧ�̯�į�����JG��B���H��92PF����8��T`��@�������alW �ѓ�/���b�H�?wJh��C��*Pkk(�3�ԓ����0&��p�l�l��R�}k��3�l�c�^�AJ ��8�#�) ר?�҂��gK��D��}���x�1�c��"$ 1��▾���[�\�9gcja��*�ts�,�����xCi�,�7�@jz�Ax�֒'h%bqZ�2>�%o]�0ME��O�حh���P�M��1�~�L �?���3jU��8��z�s7�[��|c��uw���o�(@x9,�>W�WK_�L,e�ng��nd�C�u�Ø��]��N�=(1g����YF1������}޼-��������f�*��Z�I`��m��K����{^4<V�'�
������W��1#JL[3$kX��ΰ��ZO�y$�^KYM���v��CT�9����3�
kl�a��z����*ds�ɍ=n	������X%k������b�7��"]�C������qm՝f���v�E%of�=P���K�"�e4���?;,��47�l1n��gآ*Vf�poy��cJ�hB�y�&����A�=ѣY�$l�fDS݋�u~37"������l}�oy�����-�<��wA��pyc�r���;aN{�&�J���.%�<�g�qA�r�7H#f��M{F�����@l&�I}\)��	 ��%d�v�ۭ��)Y�Zi�."~/YꩰA�w	JR5�04�VӅ.X�nB��s�$^ZsC�>�Hf=��/_�yy#�m���� �Z[U��W�ׯ��g'٘��.�Yu&�����3�	$���!*�Ƈ]��f1��Bؤ�h&��� �%_�eO���\�A]���lR'�C �[����%e�"]e��������Bv�vL��u��e����3��X:b��~��׶A����6�W��e#u*?��x̶�a�j%>�1�Tm��1h������փ^Rj3ptF0�p�}J_��>�N@�BB��w�?��+$�
������G��)����q+T�;�W^t���pr��f<\}��׉�&���ޟJ�^n����?G<�5�����)7��C[�\� v��}��� pr"@;�lJ�JyS�
 ��&Q���Rac\A�^M�U V��<��J��l?ye/K�PF��yz��I\�L�E�Z��8��°�+"*ǋb�Eм��`I�IR�P�#uI��j���1�o w��V29�ZwxڎY@�\tk]�����Sk����q㸳]����:6����!����h��CmcT�-���Tw ��!�޻+IĮ�&�ʯ�Cg�b�(�����:��V��v��V��}#��6�G�_��F�a�����ZOnK)� ��Ve�O9Bz薟��?���D9���/�z�/'��s��e�+�	 �mƉ�&z!i�i J�-<z��>�l$����/������j�X�צw��}F< �ɜ˰)k2�F[�4��hc$�H��$M��C~�dx����)L���	7q3ɏ��b�-���-G,���'��[)1����l���[�H�Q�%�񡪉94Ho���@(VP�'*�zƀU�)UQ��q ��e_�NQ�`!j҉�Q��+��3��ᔭ����\������O����XtC�������F��@Ey����ѧa>�H���v��M8�Yxi��G����n�J��x�����NB�q��$$��[=�D��n���j�9��.���,6!�%����{^>���ep��cںM�jG�v��B��ô0x}'nWH�}ͥ�yV��tn��������o�9,;�kk'�;��D>[`�!�+�9�bK���ʾ��4����0s(JE*��gQ-��� �4@�����8��cV���s<EQ���ў��3�t
��K������=R�����56u�j�]�b�u�$�</�~�J��i��Zg��a��Zc�c�(rX���w�s��W^$��(L@��|�2GN2����m̺�|Z�b��U(�K�pг����()���o��T�3*:ܦ�&<���ɄD�a����)dj���Hi����uxJ��B��T�@dT&9���Z��}���g��r;/��T��+�/��o����T1��$�-4
Go��YU�[[˾+h
g��	c)-?0}���o���<��!G z [��C���?�R��� ��L�,�j`�BTq軼iȟ*��@Y9ǁdP �����DLn4�̪2���=f(�x>2A��K��Wh�p��H�H7�M�I���� �a����v���-����'=fS>P4�N�C�)�a<�pɚ�Ke*����M6���jR/+1HX�9�k�4'�55KP��衵��vǺ���ܝ��"�9�{&�p�R�(	��HѮ�g8xtH�R������+7�.��㷍�00�����-�x�:Yd��5(�U�7*�9��+�1�R�['��(2G��΄�\ິ~��Fԑe��)�г����2cB��]w���k��>��c��*f,]�5���r�$ȁ ѱ��.m�O��T�
r�Q}Z/6Kf��1|���ba���cq��Ti� 7�|h<k9i@�7w0y�imm�Q�xM�=�~������r�L>oC��[8X�U�NR�g���J!Yw�Y���X-�[q��m���{,�D��3nWIً{�����V8�Q6�D�;D~����<簬O��r���Uӑ)�z� ��9�����y�7#B Z��rꧦ����$��9V!ui$�/�ly0�u@˂(XF�u�o�,��4s>�*F��N,k�B�un
S�]�,�`���Gu�X�?���1h��!si�]�m�Oe0��dX��2;�p�:|�CŢ��6�O7[chR`�-���T�ƍْ~�,�Q��݋Goz��X���L�����]tDO�i83��XU���2���ylJ��+�
]�9��| �,�$� �wR#Iɘ֐~)�>_�U�q��a��+{e"
�9� ��
#h�xJh��E/��������j	~_�tiD��\@�;3$%b<�}���|c���|ֱv�֟�~�\�8"W���#�=��
H���n�P|����w���$)��g2n�1g5�f�eovC,�,A�A�5�ؤ�m�}�0q�B?���Rx��=�Đ�����Ho�أDh���M|د/��r%��,0�*&$�r���� L��c�K��B��OuN��$,Ͱ&�x�ܣS4,�q{e|d���'��+�;�MD��> �(x^~���ԑ�l?��
����"Ƽ¥��<&	�	���|QH����)^r��$X�uC�� �g��=T���uc5���l9?!�XY���5����!�aUV[;GE��r��4���tU��7ԋY��T|�xK�/����٥g�L��5�3��?$cj�����%^���p:��o���o�(0���7 �.���T����.\HM�9��G��g���#��=���L9'�h�>���T0��TQD;��*��t��`��yٺЕ|Ū�Ve��H�������������r��V�ߖ��˥B�
�����Bj��k��v�
��b�
Ņ"T���)M�(�D �"�Ɔ~+����KR����0�����R��Am�k��D��F1�,D��f���C0����`�m�0n=<��Ե�j%�ݐ�4�i;�K����(²�1�
7��A�H����ྐB�&~G���n�\Bc��b�R�蕔s���$��ن���`�V���f΀��Ი��=�`�r�������)���[�uRR��묈�c�W�/$���IƊ;���	u�����]�Ň��x��������*^�AyU��)�yI��̾7�l�v4������!\�E�T�	ͳ���%=�x����M2�:��7�6�W� ���gs7}w�m	)�ؒ$_�k$�z�����g<�w0�Z#�.�x�m ��(�+8�i�cѢҫ-�b웵����i�-^pD�+* �ߞ�y��Nn{E�{���(����c�L�϶8����]�jW� ,�]W�G���}A������* ��x��ۭ��!h_��p�/r ��(��&@�b��v7ݢ�l@{2,��S
I��+c0�@	�d�&���ش�/=�[lRk<��Vh�!��?�#g�ex��и��4q���Q=��tE~A���}�(�j�l�*�����$��ja�qR�^:�+�QFW��O�O�#�^J?M��P�j2��%>Eਥ��|e�(l�_�ct��ǚ�P�d-]%}�O<3�5e�B p-�5\���T�4";:{P��"ߍ�hR�h.��"7��� �!!��!�y�ܣ�!�����C�nS����~	/���x�]����a a5
����:W�h
�����,b#WH���bZ��H}��&���
��e�Gʧ3�X'�I}2���X ��jc�$���"Xaӵ�F�6��B`�V_���r�l8i����T���N*�u�:^��BACU2�b��>�d�p����c�����k����q��?g
j��C�8~��I<���p^kG��� Dn?�M�_�^�t�Ku�����x�f���k��"0�c�cd0��3`�sr\bȐ!�����0_(l��� �(�E&���pd/�rX(��m�&�G����+zL�EɊ�.�+x��]$��b����%�,�&onb�=?8ٍT�A�)u�� Wb}&լk�� �#U*�c��d?�W���2$pi�����$;5���n�+�4�}T��c+�AP��(�<�;��q�z���+��X��F�+���3������9{�	Ň�n����@��eq��	y�3a5��%ʖ�0e��p�I�喋����8�8�y�S��_��-�	�Ћ�8˵�X{�k�;z+y�g��� �uE}i��P���G�0���Xv���z���k�i���bFE�h(3T4����bl>f#����TQ��v���	�;Om�-�w�؃�g�+���N��d��uP�J�PV���<���"MA�'L���b�K�c������#:PH,�RQkm��(!����rȍ����hq��o L���S�51Y_ث��=�W6B���ѰJ�oZ״^�O|&�'���9�@ۅ��=�d٭�qD<�$�P�qV*ۢ�:�h�-n�ܳ���pN�w]9U �Ƙ�	j���P�|��$�i� �P���	��=ie<�
c0)�A��ˌN)��
�,������l:�x�F�C��jƁ�������,;��,u�\�+n�0�>��it���dl=�X=�福9k����%A�X��Qþӿ�}���Y��nx"o�$�z�"f��[O�ُ���arٴ��!�*{�����%u؝VS�*v�P~���+��4������#�^�����-#}�(e-&�}�b�D���o����@�1�\+���7qN�٢�*�p��74���*U����u��O���#D��W�L��a�B$�i����=���#�by}��P
^%Td�=MC �kx2^�Z��?f6����8����%�%|*��ً֙��O�P�fj�4۳>Q2[���G�}8��u��c٢��%�vn�V�8x)&����6g ����)CD{�mѸ"������m�:s��nu���0��|�(��G�t��RAB�H#���]]{+��Q��Ud{!7��%�ݴN���Nk��!�ߎiۍi0m����������ulӴ��qR�iM.�Յ�ok����z���9u0� m�Y��0n�*�c?7�{6R�!Qm�Lw'�V.��/����W���������i�)r����w�'��l�X�)�I�K�w���-6:����i���9���璦�,�W�����V�$l��"RW/Bas�el��`��Z6znA0�㡒V8l��8b`��$v	���Z
��`���M�NJ�)��9��_��9ը�c؂�N%ދ�(�i�c:Ib)� ^��̄�?v��eo^�^�Z��n�H�b��%"a'r���DN��B?yo{��J�b	_/��3�R.�Y�Qq ���c��V��n�-3�/J�|Ŏ&#�4 ��o����KK}]!�r�86��]�߭FA�΢ ��c�~kv��s�M�:�]*����x��Qq��Q���/�x���je�>3�6�}Э���T�^\j���g�� ׽C˂=IV_Zl���w3q�$M�<Ƞ�T�06_8�2p�w[�5	bw�6�\F��g�_ؔ�Φ˖�T��4��v�L*��weB�zQ�@Uj"�
�~�)н�
K�V���W��C�J�پIg��2f8U��_�O��^�=��I8@Ǯ~�p���	HVk�ֲ���6�'�����[p|��nc>�/����N׬X_�ǣ�R��H��_�/c�������I�����]��b�'���gd��CGp>$p��BE,?t~u�ǩ��̫j�tdYї��dfp�A�[� `X�tLWЂR<���C�龮:6�n��F�����o<0F9}��{.�+Y^�jRj��	�C}4�"҈��Q�oءꀳyvSA3�
�y_�@����j�;Q�B+�ȱ;���ǋ+�B��]զ	����!�Pxxrݎ�5�1�J�+,������-%*�+�>�
�cq�L6�`�0dI�w`j.f��M�����A����"��!�8V�+.�����Ǒ�{��P�w>�_������0R�� d)ڊ�J����_�i������y����m��S$��d#o���bAp�:!^(��,��5�eh  ������
$pT�)���E(`��:�GZ�8�;�9҈�N@Z\Ei����J�]���}_�E�B��	(cѶp)��+��fȫ�F��y0��O�|ia���q	O0
��l�훹:hs�I
�`T�2n|�b�e#eh#�M>~i���Ҭ�54���֨w$X�n�e��.(7���W}��������A~r�p����-�)�xQ��?��S��2�c.�ϒ��*��R�I�	f�^�@���.VK��:���Q�!��4�oQ����*���������f���ʣ�P)�����@$Hb���Ȉ��u� ��/�J���������͇N��x�X\��ێ�ؖ����z��k��f� �k���.�h�=�E�'���$)^W%��d^V<�_�t���W��S^�^�Q��7�^�Y���j���쪞`��T]cN�p3����<��)=�5���\uv��P%B+p�?��DI~CP|���:Z��6,����Aq�F9�������Z�5x�ˉS�?*?`"*�Jf������J2����x����6!eT�=�T��}�
����I��]\߫! j�&`\Y�!{�|�G����a��.+0H�ǉޚeoU8��o�J9wy$AH=A���\�ɍ�{�@�Y��޺~V����4��ZM��)��1��H����J�'��R뎊O@�I߻P���F���1��CI'����A{W�q���y�g5U�gp�����چ\�y*|�2�&���z��պ���u�OQR��9���1����S��5ŧi�a�-�cO)1zrx�	B�BG�rfvUѬ>��T�_��{��D�t~Ä��Q엢�x�!s>�M_�Ȕ�VĪ/[�����ʇE��!��+n�R<��2���br�����鈦[`M],K^L��C�G�P�I��*��	},9����;JE��8y�<6����T���%F�7۬qeæ�3oBA�ӟ�م(0�H�;����`�0y�Hb�FM�].�l�8��*K�|��Yq��ca�����~�5�%a�P`��,��'�t"��N����{�V���Ip�N���!�G��2�{�m�:d)ѽ���Y���H`���/��KM�z|�t����u��m}�)�dV����ϲ�j��'�e�����JGa�;��/�'9�N�W(ԗJ9����wm�'&����w~���KTxӏC�j� �̉��9����aĕgmՎk��9,����q�}��ї�l��9r�O��~H��_?��P��<_�ܚ�[����/a�|�]z[����g�6᛭U��ԋŔ�D����8e���4ɺ����@H��l)�M��1f�f�ik�XQ({t�K�����43މ�7J�%� m��\���|7�@��8{Z�׷�Zb�(�<|.�tn�9����{�=ëք�O+�\ 
-s���|��WV�~��P&�B���{I�Ѓ�=�� ��Sj���4��Ic����Z��["�����o�1Re�5w����S&�"��R����=�45VgY�p�����R�뮭�<��v(����6�Q:��Ѩ�#��͈OZ�Ԙ��{�m��s���\�]���%�id��j ��c�։4��V����7dG�)GHA�A.�m˓���p��N�:E A��1h���JZ�y��rM�Y���%��?�{!��Vg�WLPc��C� N � �6.�ۣFR�>e��Za�a6�k*����Q�UM��g����"�&�0��M�#:�5��?�Ě^ �Q�]dE�B�iHaxX.�v���]�Ϲb?�B�[�mx��e[ю�N,��޺A+��������x���V�e�؎�
?V
b��.ıu�S��lG�q��V��	������c�iwa��.�"�@/!z��S�S�`74���Iü�l�������	HR��d�5N�D��#�3o17��,�8ԏ�c����f5�������Q,f�zL����OY1�:���a:SK<Op͔Rp��x%��m\e_�7�F��Z
�B��t[_O�z&|i�_�n3�I��<�n�#ofs�cc���C׾^^3_�7�&��4��A�}���=@�_��( !y�x͆c�#x:��`�w�&�Ө.�$B��c�	��a9;��Y�w\b��Eop���%ER��ο�a:i�+��L.G<�e�;X��6�T�%�u1��1݌���R5[�8���F
�c��� ����\o]�KC��#7<�;�7NJ��,���f14̶a����(��E��$�|�������j�@-A}��6����DW���O�gs8�N��@d{(��J�쬊�֖��t�7�!��$f#�U�%��U�]8�,{oQ�n���Z�72���@Nl辳��#�H�D���߾�j���e_&��_�Ng���V(Dt�n�w�cf�P�rv	���������ӂ�)��*7`���9%Ң#�Ü<�!=�cA����;�D�@�Y��D���
}ɥ?h�&ygd~�C��y�(�D�7��뚧��;��ɏ�]�����i@7�|s�Eճ�z�uZ��ҧ�(d�z2�������5{-�:�\Ðf��ۊ��b�H�B��I��gOr�����JC*�iGu��.�y�vS��ƀ�D=9��arǞ�s��^����
1nN?�<��~vow���sԲ}�I:C#I<��ñ�|��Ǣ�d�y^ �I.5#�<�Z���٦7���T
�?�{����]��o̰��`�-}Ώp ����>���3I����#UbO�� u�0�[G�g��K@���R�r{����8���s_~��A�M����Hŷ�G����E�>�E5m�ς�����<;�t��5�m��a�1M�Qzwڎ����������ev܆�[@�� ��d/�כSט���J�a˳@0��^�[D��|G[k�/Ƿr�4�I�.R��ת�1�w�ٴ�d#)V�;����f���� ���x�-M��~��J|܃�	�����^4[ �ag�R���b�Z��՚,���7�m|�@����k�!�7�I_����[$~k�\~%-�=�Nj�q/5R
��Il4��������6�]�t�`�I~���OY��0R{2��o5��b�ct-+M|��ϑ��Dg��F���E�^�~�I	@�Q{���v����=,NR�uʃ�I��/����u��RT5��4�ωFh!����dl�K��Lǻ<Ŷ�v�g�ً#xoY�
lZ�-�˶'�zJ2��g�	::��T*�B��i�_`�($�4�6��*O�=j��K"e���`HQ�5�D��]nõ�� ��B���a��r��Ьo�d\<L�	<�E$%*��H�����#�6\��H�*��S����O���������ZM���sb	�aiU\��7�w��-C�:	+��U��k)/�	tL��.2՝ύ�O.�$����N�wj�TwxA�rd����J�mM�-b���g���Q~������S	x�Ǩ����m>o�aMm� ��	,EФX� �39��5��W(( ���[҉;�9�H�M�ef�P������Ĭu�g��j=��u�@�a|�NO?FD==�<=$��/�S�E��Υ���Hd����}�@��q�/���s������	
-=x��
������z�@��R�W��L��� ޵B����1o�ȁAX�.�ԛ�uv��#�dFn��G �Y�̻�����;��p�&�\�2Լ
�v�������97�؍^�OQ�?/2Rv�OL7���"̧���z��.�/�7�9(
C��[��$���IHU��O���6\+�"�f�� h�D�z��~D����9-�bn��,fT�����GV��`T��#I\���Q�n��� ������a6�a�5
\}["�iӊGD�yA�c�l�o0���ٚ��
Nr�ݬ!���êߖ��7����	p�e�K%�p[�z?�	��߉ϰ�hq�xYw
���@U�̈́����eh��B=�����6����U��b�O���Bu�y���P����&e܅��X�����X6�O���a�s�`Z(��[�}=ʭ�Q�N��%���"�
S8>���0�$a���ټ�6-�UM����I�g�ML�Z�(�8��T(؈3ef&�nͧB�e�70���ԥB�3)]nz���4��9�������u7��M�k��Fq�F�����s �$�w>p��`��jm3|}Xr�����Js���߼��zy�}��=��^k���'�����ry^w���kt�zUb (��3<$�@
��>У���J�@� �V��k�m�_,�
��ۯ�I����A���=\����t��_޷W��V%ط̵�a���ݖ���l�+�z%�����ߙ���0��j\�:�#e}�Q"
]~�	��+��5�.%m���n2�"�Tz�ȟ�ב�ry2D}؋ե�{jrm��%x Br*�ђf�O�&���`��O=��C�$P��'��-4b%�8��u���J/��s�&�1�S��%V�q����I�[�ZY����R9i�n��Q�x���3�6[�+�¸���zw��i�j���KN���);�bH?��o=[��p��]qt������p�F*4�����]�XN��	��u:���(G�77Z�����	���
��%��Zj`!cP_���RbPl����|�+��`(s','&�j�O	���L����/i��djuq�j�
���J6��Fg��"H �7���2���F#	bC�T��,�����u�}TT{Q�1>O�I�d-\ny���Zyb�6n�7��c��(�����(�bj M��+�r��U:��N�|�(Mj�@H�am�a�â5�V�T@��\6����"�-���i>QvtD�gy�������\����;売׸��4�UO8���?'de����?jg���0o�f�Cj�N{(´iI-�J\�a��/.��/>A3D������/�_/&�&p%b��fX_ernׅ��*D>�#
22{y�VG��Q�28Z������&2O��<H�2!�E�8@d��	��<�kH험$�:QZ$��n�Ä�Z]��z�|�����8)�}.ij������+��F\�g�)�&nO/��Jq�,{q�cx�CF��{���f����p�6�J����<D�'3���i���\?���_E�hQYQdC���ۦ퉚��D���9c��*5�s�OLԦ�&uJ{���NS�|�$-ƥ�i@�h@���I#udw��߯q�M�P�1����7&�Q�R�#]�m��bN����%I��N
�>��������q{:t#�76H��8�����q���c@KG���J�!:��OJ��A�����fyo�CYH�-����<��7��fiT��+a%�/�<p/�Ӿ��Lfœ��蓙�������v������m�����~)@@[T�r@�gAU��ŉ��*pT���������N0F!	.�����ӳ���s!�3��׈-q�Q�F'��[�:ss|ہs��U��(��g1�?��:k���ŵr��^��ߙX
[*�p�\�A:1R;�#,�-Ηz2��X������Z���s�Q05�����c��m��j'�
}UubOng����56E�E4�X��V��s���HQ$e̹�O��.��&o��8�%|�Mj.
Nϡ�Eu^Q�.O�9{J����Ъ_`��3�0��q9=���;����Ŕ �Ϛ��	O���t���޺�y(�������E�����d���S>ǜY��mo#�y�=�='��҇*�p}����7>ϊ@L)�C�H{��̳Q�e*����L��eC��,#�����3R9=;$$t܂���s����Fʯ�-J�<����� �8dL23�A~��Wf�o0,9]���S�����Ix8�Lޏ��7�JǠ����1��2fx����&oS�O���BL
K����*�r��`z�K}si2�qrgX�U�`>�����ߵ4���Y�8q��ز�
w�="�N��Qo"���\dւ�o��"������e*��v�^ 8���T�<v���~Y"�x/Ut�k���%w~w�*x�ʗ��\ �L>F�7W|W��^�q>�������H��|��e�@)��I����!�����R��K����K�9�5����	��_4�L��G�Ջ7�3`~^�J��i`Ĺ0��K�	�H3��F�(��R����'��F�h��*���!�?\��u=c�y��U��!�c��W^W}j��5�@RH���!ފP:c.��u��)�8g"�����Eu� W��9�I RB���o��*�Z;�eP�0�M��fTK9]���WR��["%�HAT�%��2롖�`�������8����Ԥ�LL�����e�+�?��,�y�<-����]T�J��1���]r�����W+�)SC�|Ͳ���>�۱�=��D�д}�K�C���H�R a�i�����宮8�ao��VDԠ�[�'��T�*X�x���w�������ƴPCi�����Z��Hp��x�D�kJ�6�|����x��+
�!�T~F�����jKť!6��U-��C��.?��!�p翖��J�,˟��K�ј�5B���{��M�jOe��X�t�D��	Og�K>"��q�����z��^U9J���[�H��/�(B�W�'�P�ә�ILf�,aO50��]6��ѷ���NPa�Q�h���MŪl�ϗd4��\���"����R]��b��r���|�U)�z�%�5i�?N�lN
|;;!���Qc|q����w�K��f��%u���,��ר����mȫV���Xl��2�����~���	��j�>����o`���߻۹S�-�y��ߗI�v���r�7%}"�JY���P�l{0br���ݽ�3�-���d{����mk|�u��z]��P�&4�V������gy���#�l/�\AC�ٹ]��e�c��g��^�?�6v4��ܳj����������}��;�W������#֚7���z����~��g5��#;O��S 珟W�ZҪ��5���2��=>xɎ[i<��i�V�ʃ��vkE�\��]�a�NW���a7�MS[������$
Y���[��$�K���q�W���(!�݌sd�lD�Y�E#�1���[����.�l��c�{��b� �=��O�U���n���:Ո���ڪ=b���M �Y�f��vr���؇��^rx�=SE<�xpE�e� ֡��7i:��!/|7�t]��w�������Á���� �L�`�tE��r��r"�=(e�y�x����L�eZ-\��N�p�ߨe�<z\�d&P ���f�=r��N�'�M�~k�!�:zbg|&���>��u��dɨ�:���%���t�~Ѣ<ف{)��c��G�z����3r!�(w@�<���?]���E�}ǝ8�o�]����:��҆V#��HK#	�]�5�)�q2fL:�����_��g=8,zm?�C���C���X��,��3:�tR_ܘ΄W�D-TLpxE>x������آ@��|�_�"��l��ϸ�����=a��z�>�I�A��
qc�;l��.�fc��`n20�ea������n-I5�Y�[��h��5/y2%^����@��䉇��b��0���:$X�����Q;��5�;��{�����'��:���l��ZK���X�8aCk-Y���*x�֣��	/��B�E��sMx�^"��sx���]����C��ˢv��d��S�[]��u�޼f�L]��]7��<LF�;}7̬TKQ��X��C�?D "ŉƚ�?��1A`__/<�T���J��p��C�l�Qaj�hO3ףk?��v��f=l�/��#t�$�hl�wi�/�x42	dkT��
,�
p�"$֖�Ax�}����C�㺉�Ȩշ�Sv,�A3�q��E��ۊ>�zp$�N;;�	j���
�HU:	 i�����V��7�<�e����
"ߴ�Fʌn�3��Qn�1�8�SMF���g��|��S��]�4���K�,E$���+�:B�Yeඞ��P$�|;����z��t}o��{Vdg��ӷFV�`�dTZ#ܐ�ٯ_�a A���~o�q�/14n�[�az�r��6�I�C���'
�i'�?Ѿ�T�c����gp��
�DT�G,�{������饊���d?H����g�0u���Yn�[{�^`�Ⱦ�8��y���)��)�W��*�n������7�L��������B<�»��1/�S�/f+i�&)�"�����$v���W�{(!��P����Ԣ�.�FS?,F9ؚٰ-bu�_���
��g4ygKs�ݖ%����Bd��<CQ�M���j���Ii���e����+����5���Ȇ7�6U5�ݎu�҂7�N����w��&h0��F�6m��@���/���_F(�Y+�:� ����4k�]�y���-����=A7�Z5hw��X�7n�0dL�9�UM_'�u�2\�X��Ge� �i�rB�w ,I�f`�S.�V6d�Q��^��F����˝�\:'��mk���"�PMngI�#�D���+p��po����,��v־Ij���8<�w�� ��K�8>	=��j!h0��>��Ð2��¤�.&�I3��9����z?hs2a_��:�"9m,26m�71��:��m�
�d&J��\w��7d]�}U]����Kl&�4�VFj���G�d�W�}��/Q6��'�¾����Ӥ�>uR�`:FF$� �ѱ�MW�%��V
ƨ^�im�5<Ը��\��86�]py�]^߄"���v̬�n����䁞00��:cFT��9a5͚��(S'�c�� �i���۔e��vBVg81��d�4�|�F�r0Μ9B��;]i����ȷLWs�����j/�>ф<qM�)����M�Ŝ^�d�z�j�+�0��`Ǐ���QU��5���Y{�T zR�,�j�=7��G}(0�^Ձ1M�Y
��|��2h0�6�T!���<��΂Jj��G�<��`�OS�R7:�T��6DS��ei����+���50���J,��is���kDj#K������Je���G�(G00p� �
�[3��t�%�  ��J��af�ߏd���N��=�Mb���:*/r:���1#~�3�P0G�q��!-��79o�#�[�����5����CX�Y�/���!� �gو%�#8|'7���i����J���W��Kq@e�F��NO�3tIE�F�f���W��x���G��D)���<�3�������#"���`�&��y������l�yII�z�."o�A���E (8��n�@E�m���9?��_�t�xQ��ȇ����챹�X�~�_(]�]���"��͑�ʱL��o��Q��(�I��M9��pT~��|�>���=��1-�`�vcN��]�bxZϝ�0�(����v�k��hx2}�z�-=:Z2ǋ�U(�� ����-E��+�عW��&�b`�_�u��2�K�iF3jĺ��nz$j!�;�&b8�
��EהQ�s�ݒ��7Au�&��y��$A�D[c���9��T�P�i;5���n� �z#�u�s�'�/��f�S׎�.��Upg�tQ\M%�]O$���e�O��I����A�\U��~�p���?F��e,��V	�1�ijR��(�}/���Q�tm˯mjh�4s��ܤ�*����Y�t"3a��Gz���Y+���+� �^�h�xy��j)|L����L"D��f��6�=��9�eC(�/T:�i��QՏ&M�$J�P���+��(%���e�w��>�fc��s�*Ss.�x�`Z6��F6�W��>������Y���(|�F�0H�_ �$�-��tQ��'���拟(�r�.���ϣ��Q�/ǣ�� z2�D � ���˼(3\�TT0�|�ڦt��Y�ʡ�πD����,8s#�H�6/ř�T@���Z�P��@�+'GD1�����G��|,�Z^0���oLy���8�"h����&م��=n2QF�]��.��-�O�P�M"��'�OkiF_�?o��o��n�To���NS�q�ai��U+z+�����!�A���"�;�p\b�z�T*2�#�d%�[�qpdc��ok��t��&I,�������?52�G!��zh��fyg��pn�vQ�*<C�4�{9�`0�D����X.��h��nu��S�ߑ$��5G:�j�a��������~�N�7^��7>�Yb��I
bC�j�)>�5 h�<|`M��KA�n�W����S���WpU�������XE·����!�?�I�F���)�Ƕ�t	��j7���Z������qP�ۣ�8݋?�L� j4��&iKY�ɏ*�4)�n`E���}��?!��ĕp ��M5���R����u�������O	���q�O�erǒ_p@���Ii�{�ڭ�s�ʖ��B�&_Fٍ��#�a�!4S����K�5ZPk���^�����l��P�k"5����S-ڔ��k,���m�Nk-n5r�Iї��NEb��1g�3�0C:�eߍ:j'���I(��.�A�׺����cA����3<F��S��=bFz��{�P�ҵg[q�;/;���%��e1+p�1�׊o-��mħ_����̧�v�g���˽}⪫P
k�(ە$�������\gt��>����\��0`�|xf�6��5���G뙿A����'R}���9BM��n�� ^h�`�����"@��|E�،�}��Sl��,��!yDY5b�
t�-骣�$����J�%�/'���;�%v#��5O��g�Uc4��G~�t,5.���'�9��"�X�n�@�a�"���߬	��`���ɒ	P��0[���͗��j.�k��:�]=k%���X2)ʻh�y-�L�={�������kP�/����7�m�AU�H=�'	��K���_
+���Y�C�F�M}�{�hJ��tІ�#�5\6�Y�A��6����$��u��ϰ{��J�&�^�a��t����GF�F��b��R؞��S�&b�U��.~�>����d'Y�K�����
�D���~��|�,�6���I8����=P��lLܠ8�nB|������ū/UF��Ճ%�@-�{CQMG.�P�(�6��!�������]0�R�hà���N�4˚և%�ZZ��]�eq��1���'\�#W��Ak���w�t��9#�i�c�a��:�yE���+Z䣅=�X���<矋�N��bK�-��)g4+��L�-y��␖,��wq:?eW"��c*Α�%�����HM�V:�>�Tk���;<x������G��kۻr^����]����)�h�c�e�Rϫ�v���[ކ�y��,wT�~��AJ����U���&��Ӟ���@Ps���c{��K��(L�+I��QD4g^t�H����h !4�ö�-�ɹ����.⽛�K�.��U�B��,�e+A�󮃤��&Q���ck	D���fD��f�C(G��j��d�n&�:��Ȥ�?��Z�5[�Iw�VQX�jC�Jo���8��̯�)r���L�2���ͩ�F���ޢ�1�qS�Ϸ@h�=��w���_O�J��}M�W6`s�xI�;K}�P��ys�c�>2M�a�|q�����tqW�əl�{.A�]�'���Q����������A��:W\
<_4�l<�4R�`�u�14�@�%��6�C2��Ѐ����63��j�8��S1�(�L�&.�IT�_j*k%d�SJ��p�:nP㚩����;7���ME�y��U7�h���tk�!=|"ӣJ� �@޶�Gzx��j]S�QpAJRu3���a�1���+��~�(��sU��U�r��Bp9�#�i�$d��e��k���0u�L���e����j:��;������a,�Q���d��YA�Q�n氾���bW���n���������U��V�)q-Y@�⽺_�6⥌z��_��Y�J�x�0^/��#�VX!�B��=�Q���ޥ�u� �4"�Dn�IƢ�^~�����w$�n*�	^�L������޷*�F[�/˭���'�Mt\��ƀ
�cw�Hy��13��RF��kɼ�]���"@���'%J����e�Oc���1A�
e��'�ԥt�Œ��>E��/c�3bV�h�K�����E�JIl�����[���l�+���:��.t�e1�	���
��'�_�<"G��ٕB��Ze�FK�����-<�ջf@���w���� �{�wcd�t,�*A��򬱔B(i{�W�sz*S.��<��D�T��7f����Аp߮l`\���
��[ұ����o����N13`��rM��Oj�JX���4L:Yu��ti6�'�����e�+��d��>�t��g'�X��o��Ӓ��俚�j�N<'�����؄��� ]��$}㖗p��i4�scX�q�˿C��4���]~0}��}ת2&|j��{�.v�ȅ�f�t����fo!4��D��k�;�)f�D@;z��Bt��xX%xI/�x>w"�e�?��`��a�H�,q"#�y^Z�����Kv�a���f�����o��i��~Wq �&�_�)�띙r	�ZkYWd��0�@J�Yfa�Aʁ�BF���Hhr���Q#�����f+��qб��V�U���O�#����&��|�!m!��X������Fj���e���Y;u�܂�.JW;�a<�|�.�Q1�-ӥ�����>B��1�|$�胭g�HW����`�� i�>�htO��_;W"��޴I�	�I�6���f��VUC��=�q����W0��D����_�v��C�$)X�Ee�E�\ܥ����c	�g�`E��}�v���Q�L%�k�K��D�)V��	�^%
nV��`�Cq�Z�%���p\�J�o�
fIhbb@�~�9�a^�W�}��U��{k�7�<_��ղuٵ��*�z���"V%����F��=�2xak��ZK`���7�ɫ���~v*c�Quļ�Fq�R�9�w�A�G�Ikn`������5�+�(��+/���B|a?��|0Q8���'�1�˿���4�֧��/�dr&9������	S�k,E\|����^5��2��ߕ{�A���nO�	�M�B�d��w�D���V5�̟Jm�?6���L��d~?�9菨�Kힼu���"f_��L�����F�u&����'�xz���WOV�1WzF�o�X�n�%�~a���WKʧ7�kht.��򁂊t��;��]��0��:��4�iEܙ���.��p��L�r��{��h	7q�� � ��B���%(	�7������8_ȹ����F�z�i�(��kB�ÅUmuu��{������!޽:{P�:�B!O�ϡ��`M��������G���9��E��B#M�/���s=��q�b�dm|�k��{�)i�ɞ�����..����d�@��2Lal
�NUE���32u5T���:��h�a|"o��Ϛ߆��dbH[MM,3LV�<Ic�\v9�1�5��+�(��#*;�pY�kF(�.�yL�%��Eע,C��{�1�ng�p6g��6ꕎ��|��>�c�՚{]�� 	�<�^G����n~�~��P�L&�H�0���+�=�����a�	�����O�5�I�U���V�<ʇ��p�9yh���<�~�I� %tŜ�;��o�S���}Atqi�����-s�Ea-�t]��L	�96��y� �I��s���� �,�,��/B��K7��u���և����7�1Ǻ�k�{�z�=%�qn#��o�@�\����=h��Of�[��%��Rq'o>ߩ"����2
��b��<$�a9r��r�Dt쵩F{�v��"�d^�1�W �V>�Ç�ؤ��fҴ��m���<�+<T�(�%�"��G�I0 �jRE`|�#O/Wo��['�1��W�Z�x<C�!����u�2���r��懰ɗ��R�U�2�v6�3�*���ܜԵ&��)�)�w���8j�x� $$Q!�^`2_��G�;�*����j�F����g�#l�ִ3Mk�;�J�隔YP@p��_��;S��iu�DD�Ew"��o=(r�~���Ɯ'��ζ�]��B��6s���U24ntE-�\��V��p��<�#�SP��+�N�^��.��R�i�,�&��6Ak��}u��וF�4=����h��
F�5���5�����U%�'
1�}h*��s���)�d�hB��<��4��1/%L�l�@��~?�b�N�ȏ?=��p�BTh�ҸU�kG4���99A?�~97���U ���,��M+��~�q�������S�P<����ھ�^��Gk�)�J��R���(d�/��M�����v^�Tأ%������v������@�+��s�[��dA�z��kׅpUw�j�j�uMf��w�k����@���d��5\�P0��lR4�$D��vN�!l��M��^��e���ݸ{>�4��ё2�n{��ܕ�����}��&+�s);������Izti�$e�͠��\j�cYv�L[��V��,��'�{���]�LkbX|E��]^!��� *z�/w��?����+j��n��C�7�eu�����E�V�����X/��1��V�mD>����8r�Q�L��TF��Pb�x�"`*j{�=�W񸾵�@,ajҶ1��J�z$u��s��n �K�'�����|Z�6L����dܹ�=�L��jpC�H.��X�)+��4�K�ܖk!�q�� ���_O�B%�ۓ�~��C�	6R��3��� �N��[J٭o�EJp�)M;�?4�tȦ����*�u�E�lԙ��aْBcAQ_(��*��[+K}�e5���@��0�t��-���d�����ħ���?H��������].+�Ԙ~.oO�2$2_ō�U������WE��"L���c��Y�m� Ik�����/煉��EObY�JWr�������QDߝ�m3�ʅGg��Ev���)(`g-�3BK\�q�ѥ d�:�֥X��S�����۫�Ҏ��3ˈM��`w���dz6P�_f�XRȞ�J��Ol���Z�_��֮�g{!�AmV��y6W|�;_;c�L+�fwp�l�,�i���&r������(�����1�eEqJ3��f�f�������W,F�KnW	�3`�¡��i8݈���'�Eȉ�K�pH����R[�N�-ub�Bh(o&��@�,��PoJE!����i?�[E{A#tx%��Ǝ�O�Y��`px�F�w�`P4�˕�I���Ph�����t�ȥ�ݧ����~tͯu�ȑ��VKz�j�	�9H��QJ,�QD�>1^S���Ub(#m�γ��&+��U�U�%��@�P���[�(�5_��/�! �yu{�.��#h{��DC�C�(����siC�Aˢ���$�_>�6���dU�{��w��aku�f��q���$oO}kC������P����z���:T�v26�,σ��3Q�eUh���2�������.Ҟ2/ix��<��jyHd���Y
�:�v���n��h�-�K�QG{��(s�̚��f��鶩)��bn�E�!f���ia���7q����v����/�
���蕿qV���87ћ}{�7��b����X��(���'ag"�H	�)��y�@��r�=�1���0�2��f��
��ެ1X����#��v䆄���8(ь��1�N�^8 \���j�權�����)��3!x��Uޡ�mw�2"�G�C�h��Ш=H	x�
�N�^�E�cu?��� �)\�����1R�Ya��V}Q	c��N#��I���T��!�P��֢��`fE�Ab-ɤ	ͪX�a7 +	M��s�H�2ld�݄}A���#�9�n!��u�Ԇ��gK,q`i��M�O����/�$b�F3�h��P)�o'������U���2�t�6��pp ڳ�=�����Q���@��5���6++���T OR?²{ʂ���i��Г|y��qXl��F�t�	�8��Zp�RE��T��x�*�YM��`5A���5i� ���5�ܹ	n�b8P�&�-_b&o|�p�l�=|��='�؅�(�;Fի3�����n&����p�
fx����D��-��{�\���\Mj��f����{�����<�
�Y��0ZA&zSƍׂӞ�a���Ϩ�7	�&��"7�
��I������J$R+�`�@>��<�[�yW��İ꣭Ҕ��y.bGE�gz��I6�5��|���@���y]n�$��%h7�,��7�@�(!��g�ȇA�D�s�͞"0@aܪ&e pY�ـ���djo��seG֎[jH.���$���ܢ0�kl��]��z��<#�^�_
_Ƣ/.֦t�rQi�
o�{��<���V!8b=*A���n�]��,'���MY�mY#�W�����"��T\墚����Lsn���0@{��o�=��:}i�Yk���L�b��?2sq��F�:��@e���a@���Q���ǘck�d
q-©���]��$�\>��qQ�RN��n�*�.�&�껂bE��PNG�!���]f�\"A�L%Ĉ��\l��`Z�5-�/ ��l��~V,g6 ��|#n�l[�	,Ո3�(#G�{�0>�a�VR����e{,��S7�]s��xN�d��ҭX��"��%^ �"˦�L�)��n{/��hؽ���!�|�lY�]Dz�UZ�=Öw)��+ס��OڦS_��٠�c�a�7���(�R@�9te���#�����z����r)�~ĉ2؛���#�+_˘h`#.�w��ڍ�5S?S�@*;��R��iI߳z�zּ��F5��u�<qdwW�d�,(�-$����wf�7�tV���~XC��Ǫ횱�Fk���j�a�=d��h�Q��)͚�N�N����	{hj�bd��3��"�(������ɺz��T��2z��>6	j�iib����Ht�h��0�R�]M�P���~�"��r�gU�� �mAW��LAW�&�7��� ���0��oRn�^	"��3N�+��,�2)�\���_�YR-�m��I����{ \% ����I雷F�wկ�<Ӽ�௞��*"��K���َ2����%�����X���v�R!����A�U;�$o���	!���镖�~�R���2��z�aBIa�-�"�o�����pP�\�p߭�����]K��_5��<�:/�K�EA$�T�@2���u��o5��Q8���4|Ԓ6Ӟp&6�>%�OV�����5�p���!jQ�/<~ۜ��鱶a��Hs<mx{�Da�(��\�}T,���m�ZUq|�)`C��R}ʡ���62�@�32ӲGdϑ�i� gZ�8��"ح�~���P��ǻB;�}9�T/����1�6���@^AMn���)���x^/�M\oJ���ta%\�G��H6���&B2�pR�{��{���	=M���'���AC���d3{�sGj�ċ6��H5|�<�u��`'�H)��jtU�c�8B�m��VE�0�����m�nyG�p�n�� �Yw 
�������V����d9�@��Q���E�����ZO�&�,�:	��T6�.�?e�|�T�+s-��O/)0�Z���ڛ�� }�/g�ͩb���G�0�;`����;�,����t�`9���g�����/0x�`�ἂ�����&�"nAՁ$��q3��f<[��˖l�Ȏ,K�)C��N�}�$��~#*�\_(Ow�t
C�>����<Olu���_05��0��P�lmu�6�������3U&2'�{��6F#Yi������¿�p�]u�?dl�G
�Yb��E�v��,����s�S_!����ˊ��)�R�;a��Ak��k��=h�k!�P^J��6�J��I��$M�K?H��D ��h���Ӣ���G��{�l��ȊH�׫�8Lڅe��`A�u�a���Q2�Jwą́8�x|�Z"�O�nR���h[ �� %�G���wK�Ӯ�[e�^m�0�Ȟ�7(��09Qf�Ҧ�,�yv�*�oO �-v�
c�T�ܪ��.g,�
��s����D�ؚD>��h��k�^�k7�
WC���١É|;�|E�6����Na�/���?=�>sh�2����m��wi6�L�V	����us͇ȑ��T�E�aK(J�lg��[uD��p*�q�s;n)�v���ڛj���-"�]&ѫ����Xb��gpҼ��(����g�h/_Fh�r�pj(˚ν	qI�K���1��N��s,pL���S���6�;����_���|[jNX#� 5Rl�hitr�x��^X�(w]bdυ�����$��gt^P��*TA�Q� k'����f�� ����	J{�uQ(��hG�_IX|+�_���%��ֽW�iZP��Z�W�uG^Cm�g�I*#�GV� ��9�p/U)C�SS`̙1R���$L*5�q��5�/�9�"j��כcqP�����F��,=u����F��5���S�)8�����K��REӝ1�v�aEMmmYؑ^�#���%f�;��8I`���u���)�亱��6[�7�4��7���1B���n4��0��� ��:,)LV~ �$Y�]��*Q����A��Y�7qóa`��$fh��Ϯ��뮌`�?��Z�A�<��E��(�a}�f��2j�^V\5`�Be��3�wlAՎ�mD�[�H����� �AVr��UהȢ�{��fM��C	o���@9����*�
S����ċ`ڇ�zB����~���V20�:n�u���U��-f��"�R1˒M��
�A`Dpkm+������u��I���uy�n�f����e>EK��]e����Sv,��v��Y��E���!-V��H_�@��-D�G{�[)�U/Ǫ~|��>ڣ���b�4�o9��i����Ǣ�L�`�Zk��K���*м;��QyK�&��U�x4n��A ����5QR�A7b���n�)"����!��o]�;�Zk��]�ր�t��g)p���]䛴;�@pe2�)�J�k�V���!�t'�R�o��
KWz��EW�Ț~7�X����Yyy�q�m�f�Ǉ��6!��Z��`��;�?�@p��g��ճQ�F���	Ӏ;q�R(JNW?��Gk���v������k�Ҫ?�>c q���D��I�Liݎf÷J0N�ܰ&P+�c�"��9Ru����$kƺ[z�I�JΎI�5
}ׯe�S���U�>˯��5wM�P1ޑ1���V�Y,�9ZW��z�}��(����qo�џ�������$$A�Sß�8B�Q�Qǵ,����m�@l�	څ�Y�a^�汮��⯮�X��!���Aɣ*����D�Xr��� )m�+baoT�]�^��E1*^��:25Tͱ6��-�=i�x�F�I����(�}mN �+AX��_����,^1���@׿m��4�/:�����/����7)4Ӝ�{goiH����H2�g��_��b��O�>�w�ߞ�}�tn$g%���Q�WE�A�;X���Xk�q����u"�ԁ|�G�%�J0/�Oٶ��G�6�Z$}�p�7Ԏ>�����n���o\�~�CsEO����י�Ξ�Dp�6��iP͇&��ӄX�y���TD�#l�FtN7��*��,�k��n�uȤ���9t)A��-�����0AT�oϺ&�B'�|��z��#ʉ����/|i[n1�F��ʣ��~����
f{�B��*�v��Ys�@.�sY�����}ij2��CG���vڎ��@�^f���س/v�<��Vq�fI���0�E�.�xĶZ&O��m膘��=���)����@�p|�DQ�o{�G��YY8�����1:�S��(�kAWY���%o@WZQn{{�{z�=�F1G,��-[�˶�����2�<��>�^�A0˳U4Z�lbB:ۂN�Ð^��l,J�Z���q̐��Y
&�����>�2vH�(�]�H;l��u>���)<8���i-�A,Zo�&@s\� R������[����][9�xSB���1�|�n~$�Y�zs� �!�I���Kxvn��[���}1H1�a�J5��̞�y	�� k���p�B^�G����Ҿ���;�Wً�t����Q���P�r�ӂ���V��	���0y�n�Q�d��-Je!5���������LprZ&~H~�8���%l&Q�1M9U�"I�P>֜u~�EOTT���p�ck2�ļ0g��e�Y}0�t@��N��t/�oV]�R���x W����N3�nm��Pez�؃����08��9���&���7W���X�kjK�9'S�Ko��#�J�:��a�6d��V�����bR�M�_����{>i���A��n/ &\|]��z�S,!�0��h�<Dm��,_���ڪ/�x�.�R�s{�r>j�.UX��~W2ږ��@��<;O����9y�A��u7TC`P֏��}�$Y��-�T<Dwq�:]�����yz<왩�x�%�����/��e�RQ�R�u������^7{;�L0��?{��|︇{�́�E��	d� �p��b���$�NK�5�pA�<�Ka��ןQ�t��و����F�Q��jɚ���!��]� S�K7¡Ua%G�q�BW�F��Q����m{���`�Dxv���؝^G?d��4�.�jH�3P>�F���m푚�09��S���W,�x����|I^�ت5�J�׵I8��9���ԏSN%2d��L����<���������MJ)܌��k���n?�\�+0C	 �b�ų��;��X�އ܃��~�!|q�Xѡ,hl���ˇ�Jq������4�G�e�g�n^?�e��&��E����;3\��.�J
j��pi�Q���Hh
=é�J�s�I���R�h��cA�X�_�i	@O�4�Y����J�����us��#U]�~�Zآ�4�&�%Ӥ�C�7쓂��si_��Ȱm�� "�����@�\�_����Ã�Ո"���(԰��/'�_��m;��R ]�P2kg1^+�nɡ�>���y�;@Q-<�逘���&OB=�����)G��4�HcM������m<�^�S�U�,y�������8!h���g��|:��ݘ�c%ݟ�P�g#g�q�!�9��޼䇘��-V��Ֆ�-�$����J�:�>e�u�$����l[�W�8��Oژs��df���,D��L����V��h		p���?:�5������BjUNɿ�r��f
\��̜G�r�8�����Uw^s.�R�HOq�y���n"���Yg#�iN�1Q �'��m��>o�V<�4��}���}q�G�3@�=o���	8E�!�9���,yQ�N���#7�ԗ�N�c�.��#+YPݶ�~���._�3�Њ���5�_�3�9"�P�E+0n����E
hq��̟�$=F<���;�/���s[�}{��4�8������7�E��mK8�Q�bF����,�r*���2�V��Cn%������ߟ��y���.���H��q�/�)lۏ+)hej�@�0E	㕸-#&qWBѲ�F_�A��+��9?��vw�wk�%���b�I���t�Vi++x�i���rmYʷ��V/=��	�7�ް��G>���T��n�B�lVjZ����+���	1�/G��k�����t�u��x�m�����p���"��'�:0"9�����r2+�l� VǀJ���k��-���QOY��	]�i�l:H|ju1^`�uA��#��֡����y2�V|NAm�4"{v�{��z���&�&k��G���&��^0��="x��s(֩����t2�-NB��,���w�MO���>��4#Ɇ����|S��(���<�)��Ϸ�X�OH�S�:QgN�r7�]�7+JOY;k/��͖��l]��/��slk�rv^j=^����+I�'g��Ťf�OIٿ�����P�ߎ\�*�_6R�p1\O��G�,g�;�yq�'�E�l)��晣$�:bh��aK���],��A��aJ�d"(ׇ�W�+�#�{(��F")*?��(M�a�G4h}ݾ	<�+�O�C�޽_'�ed��}>)X؃%J\�6&���./�n*���es��&���{�qڭFq�|��H�6ױq�V�5Se�8����=f�[��Z�fA���p�r}(�.�x���A�rS����dT�D}�ެ�FbŎ�3�1u�U���ʭO���M���ˎs�k �`w�{ϯoU���8�41Ő�bJ�QӑP;j/4[1�mJ���`b�q�IB�-T!��62g_q���UJ��P%1�?JBf�r>̢^	+aoh�P�[?s������
������t-���?�A��n�g!��N9r]J��n���O>�aO�,+{N���%��+�:?0ǺfWSݞ=O8���r�M��{M*'���nr�U�����J"P4!GT]r���y����櫕vd/=�${���4���'rkJ����&qK����-�%m���F�}�oew��7%����|��͖��J$�k����S�7�+A�|רBD屇�g�J���!���Q�ѣp �®�3���;�����D��9,�u'�Z�>OX��;L�me�d⨟���E`67�D�H"6�t�q��Ak���ӟYq9 #� X�i�	����#�k2)��~��t�6:o���n~D�����5��|�t I-�ý�ܪw�u��Ą�˥��.���˸�"21me^?Ք'I$:��u̎xr6���ݙ��͠ݲV� 0:�~�W =X��;���&�OH�-��Y#��S&q"n{�������R3��6v����yibv ';V/9ud��z��I��TH>��e�����Dڍ6�Q;;̛�a�T�mOhr��I�D�bfZ��/5V��}/�Q�b�|�լ5!&��0'6�?3��.Q��j�I�"Pː���Ap��Os�9�����YM6���g�V�Ɛ�d߃�� �K��v�f�zN#D�ԁXO���(Y^�kv�.�������t�[��v �x�erAb�i�]<t��LƐ�u?�sjI�D�[�iϙ��(��&"jQ���#¹�5Z��̍�g���쉣�ۆ���I롁��k�9D��4���0[�����z�p��X�}�B@���Z��chu^�������ԃ���p�d�	����{]΄�����.����R��&������QR�����3e�vT�|v�����',z���z�B����+�)�r���6��3�k�j�����o��x�
���{����s�P������6A�Z���k��ݷ��٠��D�S���pS~���1�CLË�%����L�z�R�t� ���
���%R�F����2DḰ�w?.r�Z��V��!z�
ܿ����zm��&���^������YUf,&)N%�<��7l�݃j�<dl^�[��F��@oU�/y|�x�G2�'�_���a���E�		M��wB�3�~g��f+w�D*
j6�n�UJ�_�@�I&�F��=�y&aK���Q%oN۾��gU^ꋁhGr)������C(��PʪPJ���ݮj#~����X�E�����3�c��6$�ws�|^��V�:b�'�dA��á]��W��?L��*��J���-z�<�n�H��@�/�H=o��<�r�?#��y�8NLL�>h�'D$�x
*�٥��2		6#Z�O}�=D��ش9��G�{��^��qi���xAe�`��?OV*��#p+(��a�����dK8}4�K<�q�K2���� �����@�
j@D�;�+H��7Ek%܈L��� Q����+�L��/�2�q6�r� ցN}�ه3�ׯ5���z#��	��a��n���J|���?���Ip���9��!/��y�8k��C��j.�a���0�ᕒ��	�c��+D�q�V�^�^~��k�T�
�>�����z :Y��\Ȩ�.Xg3���z-Yr4F"���>Ee?c�#�a�QS �f���QR�v+�>��:�zfIH7�k��:�d7�	���fE��v�X�LC���s�,��Cw(Ĭߢ[ky�;E�*=�ƒ�9�?Qq��w͑��uЅ.e�na?���z��h,z�{����E�W�e#4M�w�H��,'c�'�����-�����]�C�&��U�K8�)�p}:l��ɬb#�\���J��U"dc�7�@n�;{�J��H��M�ƅ [�E���������AG*,�z=,x���@%����r�F5����ǣ���V8,�&*�*KU�jko?�gt~��Q�^8�����$`ة�����������Ȍ_Yڦ�w҄NRkJ��R�H��F}�(�M�V7�!���]"g�����V�ik�1�s��>N�1f����x*��=Ӈ�[U�;���R��8QM�>��b��'��@X+��<U���3pv33���Q�a��������rčgPr[z҄q���zݫ�d�Z��p�{�b-q��������~�+ʄ���:�rM���&U!Qs�:e(���_��M�Ä5�r<�#dF��r�2��\Oj��|be��[W�|+�<�O��=���@uM<Nt@lN�zp�ЊO��I�<n����?�3��:�=/�d�ng��;����gGct��×��pX*���	�ily�+���	�L�s��V�ê*A뱷����WG�>�Rf��t � b1�06fy)�1���|ܞL�v�=�#���*T�yg���������1I���޶�������c1>�F�u�`@C~z6�le_G6/Bp���@����8�إ�T	�;n�N��{o��H�8J�,�c�o�M�{�J���9�mBl������N����	E�?g�@��ܼ�:H+k#
NE���W� R���$2�T	�6eK���z�]�]�]D�l�لE�1��=n�!�o@m���u#j��I	�P�D^�t$܊A
�!���Y�0��	T��c�^�i��ґ	�?�dv�7�{@�f}�D�g#� �A��/�fֶp#P��xڕ5�5��А��N�]e�w�t��$ㅈ�ħ�Z�Hh0c�Ldd�o��7�,�f"�&$X�AG����ɀi�:�*���+N������$hRÞ�1X�ȃh����U���G����<DW��� qD����2�2 �"�`W��uiٴ.��d�^i�+���F�f���,�}%�)74�-�%ӕ&�r�)5qn��g���a�[!�^IP�<��>�y$���?F_�&��G.4��H�{	�}�08	!��ך�-x�=���y�;����V�|_����6�,Y��[!����-�1S���O���Ӷ2g�|�iS'�]46�ۑ�#&�f�
��j��n�6� ��{p��A�L�deeOZ��Xi����Z7S�,J=ĕ���v�M_�8(�/;9��Pބ����ӜJ�_��;�{�:{���5K������#�0����CW{T��������h����I���<��'o>�S�����c��e�P淔`�}M`�`fcM�|6I;�"B�����B4�+�Z�#Ka�CB�P  �f��L⮚jXxA��	���lv����/��ȱ��0~�-��JYZ4����F�R�M'#XJ���>kљdg�o��f�&�8�.���f��g ��2S�_����A���ض�䘓	��[�7�9\~9ٱ��9��kKʚʆ�+��&xC�w{���8H�%Y�H�$�V�8��0���yi@�n�A1f��7�Ӵ;�4���)�d�lX,�r|��s�OO�6���,�ۺ"Wn�!(Pb)U�TXh����f���Y�|���c3���%.��l���kZ������%�d�W<�68���~���ա\XC��zs���q�D��w��T虃S�X����X�����\���7��9-��5�=�-���H�:;{X��Y3�I��T��a�I6��_ �C�6�@;t�
ue7�v|'3h����-<TOk~ �0T���o"�Ɩ��o�Z�
��b�Uց��2�� �K�����=W��>i�ծ�EHt��߻�J��Z���xS4���Go.����0|D���a�>޵�H:`~�ū~�����ǃe�i�s�9�����A��l�����:rc�;n�6�Ȧ�la��`�sx��J�9�$ߒ	!�-��f���mbBH�B�}�u��Lt,�G$Ns��?ɍƟ���֢���A�vB%O�D+��-��(XUsM��t"�t��Og��R�~�Z���@A��ߐ�%�M�L�8�[��kT������%,�w^����
�VT�9��z3�_H�q���6�_$*?rW�tRD�1�V���,gY��pO܀H]�c(�������%��_2��(8�
�^H�k��NmR.����3����j���8��Wd(R{Ҭ_Ls�p7��[�<��»����'��֌u4G���5��M��Th�u#H����Js%���K?]ؘ{T�Rx��� !&�Q���D4�%7^NO=9|b(�iD"�r �������zxA�9�DU�Q� mrp&I+Q�Wq�4����6����#
z��lO6y�q��I�	��g_o� #e -�w�c��W�|���f>S�7��-��@����|X����l6�O���r�꙼I�{s+�V@�w���)�5��O��#�:�@x�,z�f:e������4i߅7�VL��"��"!��K�e��;����[Ȅ��LJ��ʠr's�˓�j"�r�7U��78�,���pN�yHš����[���z�6���� )a��ǶS�r���b�B��i���P��S��O�u�Q��~���g#=��-��jr��x��	8S�L�ChL)�F�5�������7�	|%!r��"k�ʃA&����14H:N�<�vu~���5@~������55Y�}2�"Gh�䧜P�RŜ2�T�bZu0�CM$�����|�ki��ڪ˄�/�,�&Zy
��3�0܃�X��1�Up� ��@ku�xm���� ��?T=WT�O���ʳ�*.ۨ0�y~Q&O�����JT��%�<��3mf�j̝`�����Jv�:_���f �j�&
���	��>sa��]PF(�LB�A����)!�'�pҌ�P$?����7�mʉ���[��y���7�*m�UMMҩ����9d�R����5��`�_n��q��>��nV� ������>Y[���J$���n������8���n(k���@��E< ��K\����*Eч�_���{4��1⃋zj���E����ٻ"r��]�����O��.B��0�oK�ݪu����P�"d.ƈӒ��;�[����>� �ރ�ɓ.E���<���1j'~ç4�}ˠ���1�z��{Ę�$v$��iűRL:����V��8�+۹�^�ײwV�l�Q��]'#��AHU��O?5�q:v�|9>ug=oEVn���C�X۶��ռ�,��Xn�\�f�&ϱYXȧ9��4�_^��;�QC�"&�s�4C1V��_��%7���T@4�)�v�C ���e���H���9G�0`�>��EC��B�]��&n7�hlm1?�(^�"3/Q��亟���r��g�'|�U�ϬѺ��������_A]�����+���^�;B�M����#�>(��
y+%��n)��Z*�l��Zٿe� O	��r�����#ϼ|�o[�[�W����'FC�����(v�uNAr����Y��L8���4�LV�{s����i��5g�,m�z���͇�^]M���-&1	�# ���5�E�a�R3�n��`��:�BZ+9��X��0���B�A���9cV6����}��mD�p�jTZ��B�D$]o�w�yk���TW(1�I/��uU�R@�N��� �u���}����y�����g�XՉ߆FN/�Bk+ᩅ�PSGS4��͉e'l��i̖|X"�����<� jĘlh�����Ku��f�dJPIt�Q+�V}�����mFxq����}�#�(��jT�zA�����E
]:����&�7sB��B�cgݗǩD�b�������FW���EP�L.x/�+�O��ZP��E>�kG�;���}&/�2�Q�7f�K �aN ��<<�JR�4�V۱Nπ�.[�c��]���'�����WLr�E���[��U�<畸ݘ�"(x�2��'��nI����p�n7�x���l
�� ̧�K{m�v�9��8��r:�s[�����:�ݑ�\��uK�<��\N0Hx�;����P��Ym}�)K�N�����]�~]�+L�5Gu�l8�rzqe�;e���3asn?2�̃4�ˢп���� �FP,�'NXb���*q|.%�
wt�������w�Zr�����˴��C�Е/	G�L�6 s�N�hns!o��2#��EkK�*���q�o����D��I�5�R��Ob�ZvI�Ij�:�&��? T��ux��&^�D��7�yE�˂\��w܀������''=s��?����A���r]�l-3�{I<]@1��Zq��H�#�M�u�i��(��5��K��aN���T˙�^�,�F�Jc;ߘ%��D����O�����
K?U��B�rjBa6T�Y܆�˪c1x��P�`	������>>:�f�7�_���	0��Or�vy�H��;�d,��̐�
�h}f�$:}��p۱@!l�nv;��z>���݂�W�b��>�/P�à��~��m��n�9΀ى���K5��q��uS_��t^N��g�� �fq���N��԰��!���ݾzK*�����d��k���K�	�1��f���Jj(�_B�o�jlo ѓnE,X����'6�i�vb��'E������v
c����Ȫ��n��;�9FRGe�1���"������xE��|��ZU��YhJ���!�L��E=�kx�C����D{�v+�h�O}�̓r� ��jC]�2����֜^��U�FV!*��Znϗ�`_aZ=�e,Fa��e;]}h3����VA��^� 24���q�!��=�CA>Ue�>t$Z���^D=<��d�bi޾��c���ed9ʯ�ؤ�> ���\C�H�C.��9���u�Ǘ�q�y+Pb!�Ҍ��[��A�5(�־o�*dC.�T�h�{,�e �H�@����Y���hj�;l�5����od��
��g[M#R���׷��w��-=�5K_�_"�|��s;��1=�����^:�0���K`�5��;䡰�IA/�Do��H����M��@�|�צ����'�X^_{[r/��ij�n����[���?�5�Ѱ��6�4������%�^i��鷒`z}ѣ-ۥF�u5�ǠC>K���;�wna��/��Xf��<�6�>?��X��i�[<{<�+B^�6�c�)p�L]���D����|��mm�v�8����{X)^cr��I��y�e��qP�T׏�rX�F�V�'o�+���/\���Z�b旋	djxE:ټ��1�gH��X���1 T_�HX!���_�����3[��H�jI�,�n����_|��o���Ғ듧L.GQʲg��a3G
� vX��p���Uឥ6�#n��{4<����zF���H>��-��*AU�/�2R����9
�oߺ��m�G�^��P{��*-r;K&���2��ІP2)I�bkn$�"�����./6N&��QV�<�:��Q��qӣ�rN�+�K�	��B}�G�Kƪ�U�FA�JNd��8�%1�~f,�`�$������U��:��N9?�sU������ ��Jc>���(�����b����?}?��@�*��z�V����C��U��LenO�i��Hc3��ٞb��ɵ��+��䶕����x��$`;��L�<?"�n�_>�P.T�(������r�;����(k�C��%T!K���O��LgkP��j�d�c���B�鬫gP��s�[���G��,4BhN��1z�8y�Mq����.%��W�W�v�k�@Ǉ�?e��4�������7��Y�yu�#�V�*w��t�ݺ�����\��*.�(kj#Ū��y��v�&��J��`��Q�'�R�����o�^t6��o$�ќ�̽��1Pzy���BN�[�"��,�
�%����!F�3�1m�5����L�O��4�)�+I�`�R�G��<�`"�s)�3�gPe�rG}	4?��O�'Q�о�w��3��8��C<%���'.�-tR�ІQ���-�_"��=���٪�u/����-3��vѧzO�љ䩇����[O�a��&{��]�Ff� � {4��אJ�o�+���%�<xAjR`��4s@��2K���0�����;B�Wi�8_S�8�-%���}A�!��x �S5��*Ge��TtDF�JG�Y�L�����웋C/��#�I��.���L)��?��י:z?�!� GH.F�
5��	nT��Dt�]h���߳]�
9�O�=��Δ���uɄ���.%j��s���VI��d�a�th`�Q��ͱ5�N7R�eN�Ƹ-�y�a<bX�@a�U��鏮�n�Kuȵ6�e�SK1s&a��e�q�n498��+!��mqǥ��sɞUl��Y�����j��J&ތ���&B��#c?�Ęt�z0�g�rF-D"�����~H���j��M���`.��v����}��g`���uw:�*�)�f�9eƸ����o}^�<���,Y�4zP�t���7��������+3q�bS�I�_�"��mxTFz�B՗�^Z���kj3^Z�3��B#t)��ck����������l�!����n.]�1�7�G==C(�ҵ9g],2E��ٍ�Ʈn`�����){;�y`��8m�Qf�NJ��,�2�2�)�V3�I���>�G��}��7|@����$�B�퀺�_��rM�=V��r5C�H9!V��rŔ�z.ͨ�&���C��~�l�_��Ɗon�o+�%�,�4g��Y@'<,�9J���}��>T���(P��<�o±�P
y՛i��FJ�u'����,W�q�����ts����ud�濿�9��Gb���~D�z@63n��F>�r����i��o�Z����EK�(����-�G���QCh�6hY�AOא-Q��=�K�A�)��jo��M�m�e��҄�%�'̟H�#�[.⍽��*׈�b��D�P��5��#`��w�^����%�(^�{ؽJpK�Dm�
h�4���\�?|_ϑ�l	,�gx���ڋ�ĺ��D®��$>��.�S�%�d~H� ϩ���� *Q�p��x��B��r���&5��R��Ȥ�}��[ï�}�"�YC��Nei�kf�n���eMB��3���7 �Q�t�j�C��3+���/T���S�(�Ho%P�Mb�C/9Kt���]��-_���xJ2y�ܰ����f��J\�/@I/i䪌��%��SV}pAb���9U��y�G�T��P�oNt"��SXa%��R���g�V�õ&� �j� ���-JD�6�$8��Ė}�.�t�"�AP?���Wc ��ߑgw�
aL��Xs
F��|/�~�E��yX�d����/q�$����S��Qx����tw�H�i��v~!H���|s�TP=�b�#�WBU�?�X���i�e9���I���r�1ޒ��QC�\�1L +�f�d�H�����d�q6��U�g�D���?*��폟�e�^o�|�̖�	�뒴���6|�c���FV���
�+6��~�u��S�Ifφ&��I�u�v�1V��-M���ͽ̭�
\� �}��1�|LU�������>�a����C�R����)/H���cWs�1����I'���t5�!,����h*ӳs��x��vH��N�r�?�%7�]
��
"�D��V�>nL�US�B���9�i���,��x��N��L�����x�ŀhJ�c���E6㑽�+ ��5�߷u����3���j�$������n��=y�#��X�{E�o�I��3�M*���s�Ӥ��1��i	9�T�Ӽ1�u	ק�9tYw��N��U��qТ�.�C˿���A�9z0�ᮽ]ђɿ�X�>�j�V�W}=/������+ŭӁeB��}G)�����Y�W�D����d-Q7�mӮ ӣK�*�ߩ�[歶C�$˵��d�硞10h���}��M���H��	�M&�$�=�^5H�it�=�?#98���!�6��<ܖ�����X�0��MNc%�H|:2�&}ӹځp�������Èww�k�I��
F�X�y��@V�[&��H���U��/��p׵������j��u��B��v1r�?r�_M�Iީ�����C� �]��!<��8����9�s\�Ь��!V��+s2���E�K�{ݭpzЧ�n�y>.�x�"+M�vr���i�P��,����l(~��lKAA�`�P�E��r�d!B�h�GPG�Je����u�
�VN�;��>2a�[��_�ߙdN��.|û�Xol�w�,��_�,k�N�G��.41b��k	���Ŗj"�}�pM��S���Ԕ~�t��/�G��ߜH���j�0!-h��Bru�w��{��?���iT��=�v����~ϔ䜒pw�W_�IBdl4x�̐�g�$s��K����8���.��K��}񋤑�8a����M�B�=�^z��p%Q���q�:c��i[��'��MG�Z�ǳf�㍘�e��yL�V~�xpO��ǋ �"q���/�Q?M�m�v2���!T�6�9 ����O���� �#e�	dv4:樁*>!�wd�����ԭ)K8 ��W�D����3a��@�����-�S�wj,�'�K$�rf���rLj��R�@�����Ի�K�:��w�.%���E��'%Z�=7/�Veat�czm��#8����Pp%� ͞�B18h��H�G��W��#�3{C�20kA���o�;�)k~ׅ�e�e5;��2JB>�.r	��<y�,"����'d�<��v���Q|^r�'N�uH
o	������s�y�_�C|k���p�r�G�R��k�G���m����H��t������\�B԰Dx��s����h�vr�ӶM�J ^����3��DB�q.��GF�Q��e�,��'L�e�83����ƓD�5k�C
<���j�fRXg��}_Sٶ VQU�c�>�Մu��.���7�&M�5sn��so)l�J�P�kZ}�0Y�93"|�l�U�(��g�|u��m�Zjq�Ѱ�9�z�4g����Ǫɝ����6��r����^��_�®�y����@�Pܢ�9Y7�Fx��i0�6��p�6���������ا��o���f���Qw4
ڼ���H�8eq<O}bS	�y�+�!=Z��>�_M;��iw$�T�)�r�K�/!Z@�U߱��7�rG��$I��H�[g�>XY��H�˃��g.���)p���^5c�Ԇ���OR����锹��=T�2���W�"{xfʕT���+����l�� �V�OI �$`��>}��|:���]S�Fg���DS일a�y�bP��̌�V2���i�N��Go���g���R����y��%4���VZ��.U'�T���pum�1S���u\ټ!$��7�a[��Y��E<�.W�.{���_�R�i�vK�H���Tҗ���w�Ѫ8�v/߂W����q��c��N��*7�N�|�5~e���c�X�i=�*V������o��!� ?Vp����}��hMv�P0�v�Br���� �?��]��L	��Q,�tv�:�a*4%%�W�1�M�*�-v� �.�ˌya��pT�I�(��E�Y�E���Qᛵԥ=mӦ��>�d�[���w�㤧>��6�(�����k�7}Z��w�Zz�Q%L���f�ۆ`[�����>!�	a�Hʜ�f?&���LB{6����|h��R��	����X����ɗ�6��o���:�I�)a��"$!��.%��o�� �����h���V��֡���NW�ѕ�9-�T 9�:�����Ab�o���i)'�v��B�o}��ۯ7�}�,�ܭ����~l��y�ЗZ�z���J%����^��	�`J�iG�ڕS���E�GzZN5������S���L�D�(����;7t��[�]�N��t�IG:Z�IB����H�c.P��γ��s�^)��>�ý$OF�c������}k %����h���D���i��f6K�zV,-4��c�$p0�{�ۛ*p+��K(�G��w�d/�0_�J�"��o���'���n�\�+�BB'�R/i��ϡD��i�`��~3�Y\HD܌��5��C��s����tQ܌��+}Z��&�`�"ա��c-
+ILs��;{��mhR7e�$c�t+��d\�<��{�+�}��e���}�B�T�uH�3&�K��*AѬ�i�<oK�fO�����JS��C��P96{�+�5�B�UQ�"��%���s7��Wƚ��ZS�ޓ<�G�u��t����:mГ �C,&e�bl��:�я��ֽ���ņ��JX9gƉ��6�3X���'��[EH�_rⵦ��������h��ٝ�#�.Rɉ�Om�٬LO������u(3�*��|�'�L��l��:eJn��L��]�ǜҷ^����T^��m[�%A(��{���(EE�y�$~^������ʇ��Q��^y �|�]���8C��f�F%2�r]\=;��ہ�r�2����(< #���٠�!�,�˾��V���f��_�B��N
�xcO��<�#�HI�@�}�n�u���$��H204TC�b\����،��\#0�+��{��J�d���ZA�-������9 +p�C���T̃���h�
�t|N��"�q�v�<��_�g�
�����"RaNq-k��L#a7�5̗E��)i����H8��:C{;ݑ@��;��f����O���P�7T+1b<�W��}Q��ƿcئ��m�� ��Ƥ��>��V��G<�#t�A��K��qG��M�&iB����"���YQ}�bU��W�B�EX��5��x���@_��K�ž�}�DD�-ߧ}��Z�T�Z���������4sWt���N�w@�t(m+]�"u_��g:�/`T�DE�)��E�dt����<��!��6x���E��`�[�p|KD�}����5 6�M��z�`N�95�7���(��ԸI�zwwX��/��`�dum}�gPD���@����h��EK5b���pMW
-��cDr�0�Tv�6��/!���>AjT�=�+ʼ����R#RLK���@��(��r�F�+!5OhT����lL��Qd�[F���V�(��y<1>���wju1Y�9�75ڸ��I�R_���8��FL��|n���ؿN���+��Ԟ	���~�7�ߞ9l��S#��%,K3t|���Q68|5IF�xQ5ӎ �ɉ�R]��;��z�z�J���S4�-���֢�G�嘲JgE<z�&:�-Q�Ϧ�.�I����<�%tNI`�J`�$�Q3����H7V=i	6�t���T`	�����:����cGx�h�"��͛԰���)��}�4Y�r?�ˮ�`7�LgT]~H���G̥�[�>L�#�cX`���L'��M�����FC'�h?��Y�	vCϫy����֊
g�+`�A*[���̢��f��Aɳzm����lzOy�:5��/�G�;������R��eB9��xQw��	�x?����S��Iz'��E�+�=	|���1Z���89S؅%@��#�`�ugs��$��:��̆��Z	"�[kXFU��e��� QX����V���:�a�; �,1�XЬ�+�zB��R�dв!� E��u�����I�j��i�0����I��,�7��2ҷ���1��\�������P����g@�FP!9���*J��A���4y�S��|x����_�����yK��ެ�]\$4��\:V����O�HD0�1�!�0&N����.����!�4B!>�ɍ�8m���x������n���v.B�n1֊��p�E�w#���o�̴D�g�l��7O� ;hGKHcI��4�p��w��&C},Þj1+��$_�ڦ�c�O�F5Z�޼7�c$`����Lv��Pl�K�g��F���w�I����T�7<K��,��N�����'d%�GW���	cɍc���m�=8���O�|tݲ/g��`�u�ׄt�n�=�!q�q��a�y�8M�s�X�r��^���#���4��z�:r�gO*Aj�f�� �W����$s�hA��˝c��(�������3�
��:`�z�Xj�ԍo���,0�q�#�?�@�sZo�f�+W� ӥ-x=�Uν�wQQ�V�h�.3\8�J��Q9�V�̽���hk�Hr���L�,��������W��Q:�y/��^�v��a�6���6<�ײw�'�%�x��\_O ��׮y�$����kj1K��*J�Y��ç��j�!:�(�W��I�Ǧ�f�3y$�](�O��H6�UB(���&n�8�R.*��l��2}�Abʶ��YP���W��$�K(F菱�}[�x�\�P
y�4Ԁ$�ds�j�wk�{��3�~���ҶK@�w��&8��%Y�6��(���~����I6)\�$��|=h vJ��OyQ�>�X�������"�^i1�IBh-xHU���=���-b`pR)�����Oa��-�h����d�l|`��ܸ�{׷fò[m�4��Ə�1��S&C���V ��к�������Q�yj��Q��"��爲�{_���+�Η	�f�9@HXȎ�r����E�Qwȗ�<G�a�?@kw-�~_ ��uĲqtY/���)Nm��&vjo6Q=�^nmVf�XII��Wr�<�4G���aRe���z+�m%O� Խ|@q�Ѐ�j��+T�S�c�g�x�c�����pH$z!�Ӧc�!�+��Z^�X�l5Z���J{���K�*ȣvA�F�۔�.�b��m��}�Z���<�?��J��B	.91�e�i��Ϋg��*�%����h��'���c���[D��H��r�7��a�b�� �,k��<Y4�K+�\��U��i#���"�z��_�
Đ�q,]�;?��`�����gx��s��b{y�[�u��S�"W?����e�Ƿ��h�L���Ԣ�)�:� ƃ��O^E�jA���V@A3Q��Hn��|oۃ-��!י�Q�E:�D~a@E����dQi�lٝL����bM�.Y���,���$���a��b���KC�"�&�xf�L 4[��vD��w��d�ɬ7]6o���t7=b�D6u)'�4��(,|v��[�9����������ɇk*�;��Y2� ��_t�������8��_"*&��aǔ�$�^m�t��n�R!TF�}?7qF�5�`��lq=8Olc�^S:�R3�)+Z���涌�"� v�IQ[i	��6ވ�\]����LR�3�0�r�5m�1�{�7i���ܝL���2>7�=X}7k9;�W�S��Qzh
�N;e�����4�t�� ԜB�_8���W������M�r�d�R�6�*�����?�-�2���F1N�!Y�#R��V+�����6ŋ��ڀS@gt�R`K��{����2���8G��ZB�T�{1%ww	�c�?�T#Hs����<!�elzƎ�3�B�a�¡�fR��y��ZN&�cb�6���10ⴠ1';�D0��l�B?�����e�����oX�sU�&����<�G����5� U�C�\��-�\�@�q�q��"��	^1FJ&=�8枤�����BՎ�H4�'�{
5��$��ʚ} �t���By�pe>��?䀷d�W2���\&Oo�y��y��DE���k�z},w9�7.��]A$ŀ
\H�ʐ��]�扥5+�O����H�A"/%��)K9��)��ӆ��6��Y��jX{�y;[�wI�q�x=��5�,�%p����Q�;y�>M�x���|L���3���ב7u
�3�^W�_�4�2��6�x��ט��SPZ8�äC���aI��j��S��8�Y���d��PYrC̄�I4͸�'~�@!�����#S�B��]X��9>xk���6��s��6Y�s�߳�D�S?��T���&��EV����Qas2�!�����5L9�B�9�OҚ�	���Ji�F4&���TI�B��������H5���v�(��!c
��	�u�0e������_zHc�S����a���J�`�*-}�(����Z�L�	���(��/�ި�#�L�e��r6H�����\G���̓@F���`���cNl�;��0�ڌ���^�ԁ.�G=�	6�_�BI�o�@�=��e�*Ɯs�iqZS�_�Í���d�TGz�bt��$z\zKiT�Ys(4P\�l��ɷdv�̦Y��Ny;��.��<p�E��1�#�8�a��:�P�7q�ў^ZI�?��T�9��M��S�Wn| *]kp�M��Rj�`�����e^��(�a���	�"������oli�󩔰�*�L�y��a��4|m�2K�Fl�m��P���gPf*��X`_�57��mP#��_+�1v����2\l�ږ��u���x��dyC!D��j_W�4CBE�E�H�N��z��Q�+��0`њ/#�˪F5&����7��,gN�eVUe��ze{g����0����@6���,��`f�ͼ�OKov��_}�K��n��:��Y	/�����,W��V�{�\<��}a�@P��+?,v�J��8~_���ȃb��|�����m�T��+{�E(@�K9슗z�2���aq����{�__����"ä:?H�Iz���9,�Y���uM����&K`݄���Z ���i�L==�P��B���@��c�o)
�@ǆ�ʛ��"�s
�b )���^D��v���&6k�V�a�]��k�1��2�����/`̰YĩI0�7�*/K5�L�M9 C�w�v�X�,��`�� �����A/H8����(9&�q����yK�'� ��&��p�Nw�p����B��jKqat�|��H�gҲ����Z��u�e���N0[d��(��{韬����H�1�I���`�KD��j(FQ�g
��`��@_/>Oj�s
�$�0D�"�>I��v��r��<��q�WK���k��h-L���3e�]�b�eh��-�KZ�)#�<�['�kwm�|�Bl.u9J�ȸN�)�T�_D9�C=��k�~8�&�ф�C_u�Ԇ.�S
6v^3�����fS�Bp�U3D�/���)mG���O3j:����eg���桌N*���[U`����8�s���-���O-�^�9W �/�L��Lm���4��PAGt��9C��ۻ�Q���R3��1�}b��T�)��/i����;`��>�FT�e�j�j�[B������Q�J��j���ߑ)�#ٮ�S"�d߯C.�)ѹǈuؒ~�� �� �tq�r���6���>uw�mԅ�P��T�fi��q��'
0԰P�DW%�32&L8 eѢǵ�<L�%�X�����*F�":-1��hH��(9����5�QG�c�-9�O䬍�Ũ���h���xbN�~�*@��r��PfG����s���1:?�tve[;�Y��#�jU7@x@z4K�,+Q��
�OA�K����w�i>_�Ê5ΒT�0����AD���(���x�#�����+�f�h�î��	u&��6�� ��|��0�^[�5ǽx!�Ս��j>"�t�J^��ό��m���0Iy�=K$m�s�ƾ�	E%d�p��%���0�O�P)�92��)�A7~�k^�рx����;9�9� ��������(k�@��ja^�z�����T7��WI�e���u�y�IS���T��H�ڜhXu�iCFlq5ߞp����p����Κ6��޼b���B��,r��5��A�7�}|�B�Oe�޷�e8���;Q��q��o�Xx���Z��t���K�&+��I��D�7��~Q�v�甐�Ʒ1qk��JQ��C���H扶B>�h�q/L!H���{��΄<��Rj��*&�E��#�,��P&�ȑN�Di_0+����b�qu���	Xl8� ���=m��:���7�]vo��$��c�pMmޏ�b$����k�aRcJ���m?�Z��RQ�� �Z��f\J-O5�A��b[bw����\?���z��� ۲�\��@\G�³�er���#�m��g��i���9�m%2�YߺU�d'(`ZUd5&ͽ]���	y��j����jMn9���s�xɈw�ym�é�����A��;�Bי��,�麾���p��bձ%st��%��y����e�����JY�US)K���N*��*�A*P&<��tdb��10{qjɽ���=����+�
FK�@*�"�>*��*��Y�����'�A;%Yα0Yn)zv����tϏ���b ��ѸL�k��̭���Gܬ�|݋[$x�mK����;)����G�N]l2���Ƽ��ۻP����#v�#�S[\@�d!̟��m�v_��>!�̕��9��
�|���OC��~�}���|
s�E@�Mb7,j�?��W.��U�=�Rg���R6��2��/(mBl�<R�8`�������v��l_���q"+}nW�{3�-���o�t��k��;y�}���{�`�����5D�Nm�2L}�Ku�cQY7�q���X�Z��~_����}M/(�� �	���z^SS�+ǒ#��e����؀�+��К껂�A9��
MGJ�
J��!A8��͠��"��dZBY�O]^���-�X&Y��?4�=H6�-*�a����=�k֏�����p��˞]o�2�&#nǀ�_���=�F���C�B�F#�N��L+����WA�.{M�$�U��/����d�&q��������aъe�r���P�;��._FЛG�)ۡzm�.��;�����Pg��h�#����?��7BYq�'�����'�ަT'W�m����Z�:�/d9	����X�t80���B~㷳������D�~X h�r�c�{�.��<"�)���Ktu�P .X��j(�:p=։�`x:�sE̬N!2N̑��������4�VxS�J�
�n)Ⱦ_�BB�h:H�J-'�������*�Ha[���w��.B��,� �����y��7�I�y-��ۀ�»�J��,)t��4�r�ok!PEp�Irk:��ܣ$_=� ,�fl7���7_CB4pl�iiH5`B[��Ztʫd �Yc��R�ī��M"/���S~&x�<�D��,�QO����>7�[-�w����g���ha�4���X�-~��6��v��ur���y�qUN��/À�JT+{;V���E�L�KO�Mx�N�L9�M�}J<^���(2��[���T�;��uց�h8�9���� ����H)W��`��  ܽ)W=�yڬvٍ�,�/W?�Y}m�ɯ�[Kg����~�sm���ۡ�b�gf�v�-�a�(>t��L
s��ٚ�h�bb��Q����ͺ$�:��=�����M�L��k�Bf���������13�ɖ���?�,�HS��	���������c�Ѱ�"/�l1����F�PX�Mj�GY�����~�R����&m��E� ���I�tP��3L�85�������O�B���t.���н	GZ$$�.�T�s����5�׭��3,�]lܞ�4������=a�`�<F;H�"�~�[��U���[��(��B[g�k���	ꋋ�/)L�M���?tG�X�ߊH���%;	Emm��Z���}L�������G�3N�0`T.g��$KJѥ�;:a��:�^��Cf��^CJd�+�Ot~2Ex�l�i�U��iZz���m�É�G��&��'R7�Ծ��>�K-p�?�����~�ң�ڒ��.�����R]��J�,C��UT>{�Tw	����=�u�ݬ��È���ֻQ��w9��ޮ&�� ��3C��8���q���;��9�\'���d��/�A���v|�g5P
ȐB[b�v�](%��� ܜ����x�Kx��q��T�(�p���vH��4�-��Նxi:��z�k���yy#t� cş�ɞv�K�5(����gs���v����-b���@Ds��M<h��<;���DP��j�޽�g��rIT��"�m�ܗ�F[f�� �������s9 =�c����cLrP����Đ�\L�b�S��M9���ғ8���5S�۹��#�9o�+դO؋���.le���E����\`�BP�SL�N�i�ӆ�(?w�X�����]�   Yƻ�TV��ɨ����x�+�Lh�7	�9q�pHz�����3n�-������V̶BM���u��w�G^I˄�pܚ$
zՀ�g��$��PY*㎙ ��� D�ң.aԲ�ro��S�q�O��-�Q��������v6����U#��S�9��\[�L	s��( R�Ò�����C�.fj�&��%e5�j�_vO{:+�K���tfl��P^j�xyr�Vu�ҭ�����%�M������&)J_ˢa��nq_(�!�s+�O��c$��ו���{
��@,ts>o�a=�&fl:�,��`^J���i�I��u$brA�e�!a���.G�ǈ+F�o1Et�	��R�Q�zx�.Quv�Ǹ�[{�[1���]tf��!��䘯��@�fo]�N��P�?A{��0��܇���_���7�r|RDƵJpQB5�S7��?I�y�ֳfEM�f�#�@>�3�F��ze��^�&�䳫��|OE9.�~4��(����fͽ_fi¬��uq�����4��D>�r�7����Q�#H����Y��|�u�e!T�G��H-�"�ey���j�(�R��$�c��~��M�l *rǙ�0���m4^=>L� �[x��1m���ʠ$k1j�L��hX�MO���om��#���\0�Ԇ��[y_TaK��|��su��D�yf�����SD�Bp���﬋��R�p�^&*�"�@�x��X
F~�]��T��ީ}�ꩠ���x���}�H<���hly)9�B�hil�<���_�uW���E�'���AE��ds`<a�b������=�����
����bۄ�. d����V���
%M�X�Y�[�|&��z�t촑�I��'�i����
:2v�O  [p���뎫>��kG�+gF%��g+�X�Ld��:�κ�XD�S�xz��A|���7�������,��f���۾}߻��
�ZiUR��(Xh� ��<	��Wg�n�*�m��5���
����*����a�$rw���B��l��ӿ^��v5�W��p�n���⥝pX�+ր^�f4h������3��b����!S;���X4��m)��S��X@u��1���a!\���N,d�0[���C���k,��@��:��`�{Ʌʩ�7"�2�XN�?MW�?a]!���_0�Iq�MT�7w&,��9ƜC��9��57��K���߆�w��z��d!�
�e0@�g�1�xrse�C�����gѦ
��V���6�
h�a��B� �8N1���3Q����.7���,Y�
b��|K_dIIu#�I�H�2�?b�̃S$\ݢ�״�Ū0ɘ���"#hc��9bƽp��G4[�֔��{�� +6@}���K+��`g,,F�@�7��d��±�e �DH3ئ�o��dh|�P�x6�Wh����։bbZ��{���IGD�*��p\p�c�ڸ �BH/� ;T1��F����WJ#-����T�$h4�n����2�@#�b�P�I�zRt5OJe�����:n�#�z�2�L�>�����(F6MC�n�	�����kx�*��3mF�����Kw�+	�y�w ugk�� ��M�F_�jK�jV�/�b��ޞ��t|��.j�w�fyH�\��|)����I�Rt��"V��D�=�+��a7i���#ӥ���P�V?��g����d�)�
��W�s�S��������`_<\���_q��T�*���<M���h�dE�_�9�A���wT�g���a��k�C�|�yk���+�E۷[�Em'`�@�<9�ُv�8�%����[e�j�'~R�g:�pDb�k����>��7U��)�I���>K:*�vH�e��C]hUAv������)Ɔ���s��%�#� �Le����*;�]f;zg�e�����^'Q>�!�����T� ���1+{����W�!l���e�CDm�`H�Pj'���\�mO�7�$A	T	��6l��Fj�������?՗�P�La�(�O�P��u�tlH7,��+�v��h��U0f{6h�2�=2��ȣ|����e��m��]�׬CGD2����M!�0̎L�w8엠^1����b��e��@�b(W�ƘU���qʖ rR2�w���aB4>B4P�`���!��/�.��]wMr����v�%e�*Bn\U�O��+�;�[s��f����z�����!��>cd�y�g����?� �&0�g�7;���@�4��G�3����|Ű��F8�t�a�Z5y^����g<�x��m��Tg�CD��k56��q�4C��b0y��5^�mO����GU�0j���I*����|�R@'�I�)�Q�o��u܈����`�6���'f��$��t)�DA捤d��4/��O�c��@�'�Z���`!lΩ�f��$W����X؆�	-�gΩ=F��b<�yԪ�tI�q���NΘ�����C[�D�T�j�eBlELW�N{�8�NbH3�ݍ���yoZ�v�}u�q�k	�v`��"�jlA��-�D��"*rk;?9�G!.OB�)�k���9��|�)��+_�&+�|�:
2���|�����9n���uޡ�I�"�`�y�A>�����)d=�������/o)�n�`����W���H'E�Ts�3��Uk���p�O��C472��|�pC�v:#�lI��;�>�������D;0����T��0����џfI��t���Yy�� �ڱ9-�����W��A�M�k��_g���S2�2���&�P�ϊ]|)JOw7��F=��������|x?�2fMA��h���,�D�*e�c��
��=���W单g�����23��������@y��fcO��YJ;7k�$k�-���Фg��e0��p�s��gp�+���8�{
Q>t�8��,jK��r��/bo�B-�|�B5ó��#u� Gh����� b14+�N\ͽ�wR����a�}h8��}��T�g�^r�s��1LA
�s��Gj!C�/p ���ڎ}�+�Ϭm��F&�ȟH)4=[�;wdt����犻s|x����13�&���y"�`!�|ʵ�q�FqE�7�
�G�}���J���5\��&AhYx�����Ae�>߄7�n��e�<�7���/��W���-�ź#t�C�QmF��B�T��dҫD�H
��N�w�}x�3RnrPp��u�%:m#��u�Zm8����7��0be�UP e5����'���u4٭��O;�m�f�qr���.���}��ݥG����%���j\�x�i�N5�JNo�ΩL�#�ϘJn���C�>'"<�P��[בL��IKt��7�/]XlN���Y�]J�C��*w���v{�>}�8���Q�FCn�,�A�׾�Hb1�]e��B4]5��VSO�a|0w��V�K7s�1�R���k8#��}���o�~޸�/cn�;���d�A��qB+��Oa��������c�j-a�b��l2ӄ.í�Q���>����~a����sS�b�d��
Y8S��Q{��� S�����۳�5
���j62��'��>`B����,�șN�Q$C��;��T�r�{|���k7���Z�� aY
��O���M8�^��{ɕDӷ��2�^܎�,�OFHkV8��\H��"�p2:�8��K�fLcD_J��RS��-������~k��k$v�JR\v�M~�-����p���簈{H@�p��׊�t||Ӆ���D|���9�٧�"]#N�QS3�Q�޹R9< ��E��E��7
��Q��{*�I+�I�Y�/��'Ec�?�'���}���1�'����m_�ߥ����R7?������6xd1N��rĩO�^Yc
{�Ze֜x�4䗠����{��u�y`��-����/>��E;�?#P�����`n�t#���m+����.�j�b.�A#\���B��hZj�ڹ${���QvU���G]��-��:��z�@nG &^�����RM��Aǘ�>~�ƿ�6��W�9&� ޤ|�Lfm��ϙ�PZc�<�� �c�Q��Uؤ�l��W��6���1]%�0�ܫr�w0���C���:����W���4-wȵ<������J.H&��U��,���a�ѧI��Ι�I�b�bK�uVj���*,�)J��X���N�}D��ޥ�2V����u�0���܅��mhŽv��u�Lw�8%�"!YV'�."(����	7E�NL\�26��X@5W���Ͱ#?n*��A�;G����%���R��d�}���x�$���"^�H�H���2���|@��ف���	hV@$���2�"]�7�I�pI�ɷ�������!S�%�
B1�*P�fb��=�>t�p:��:F��K�)c�g����D�m럡�5�!^%n-t���}�.�	ywr��4HY�F,H���ﯽ|�EJ�+�
����dP(Y�[e:.���n�P��J�3�I�Jr r�����uӳ��nt�>�����c��gr�܅��XW���JW��MNJ�b�@�8��G�:���	���/ԃ~�l𓫾��Cy����Tm��'=���+����0NN��b[��qc2�m`��
�B�.��6��yC��`ѝkzGI��>�#�^ꪆ��+c�T�V/l�x��뾌�Ts˅��^��}��`I?9��IJ�~#�H�롃/\r{�|��c.�}ov�F`V\4n��3���T)ɰ/�;����Qoc�k_�n$u5y�[��|5C�&�Q0.^3�賊������SSz�\��������.��W����SM�c������1&�,$��kӃ��j�a;�G3�Ι��/������輰S?P�):�Łx�f&�
K�"�w�����r+�.m��5{����ԉ���q�ї�yI*��"[l�/Ϭ�AMC��X �7i�<e�J�}����G]�H��Ё�|�/�b�S*���L���V�{&V�����?�6,F�����z�~*_��}#W��ó��-� .1�k� �m"	8��r�pf���9�|Sy��˻�K���<4Lk���wXՑ��*.�З���$m$������`��
�5`������/%������O���g~��A�rY���Ӄ��x��&�?��i7~��}�b�1(�36G�7[�`ucS��e�q���)_���B�y�F� e�46�*�I�p��(�r��ϱL<;����)����]��dy�>�tL�����_��k��tX��S�JS�ZE����u��؄(��;='���.8�ii��pl�n�v�X,X.CEL�j?甊�L���;#m�ֶ�Z����]� �KL��1�Rrqx{Ÿ����W�v�-k%�J����5��Uw8wd���f�O(�B_%K>�I�m��"�,����7�̥E3l��9ugy�]OΆ�z��%t{rN�;"�L	h�(��h��|�x'�^�%����X�֐�<A��u���XŌ���.g]]���	�u�V/�O�66�D���o���m!���pN)F������c�ov]���`rp���Ƈ���)�`����L���7��F�s�����#ؑ�S�8�Nz�o/�sR���T|�p����W_��`�����o���}����b�s�B��M�Htu6?�k�+�no���J_̡��j��G�D@mc���E x�1� �,n�AS,����u}��p;���Ջ�lь���S)M��I��b�VvU���gU8h����|,�r�^������(�_p����yu��b��}{�#��Y�< *��o�������1�};��<�))ú!�UBr��[�)��;�z��������vg�ߒ�	\�(��ƹ.�eq�=RUF&��{F���l��6�:m#\�6��b�rn�H��pJO�`�&>5�a��&�\�ֳ�y����8����֓����|�N!��Z��LTۣ��ϡ��bv@<lO8�^xŻ��/�vg�:��ԗ_��N�]N�.�y�~�Â�z�J"���9�-ۢ����Jy[�>�ݏ��~	4��.x��A�h\6K�q��l9��\A�Sq�U��JcѬi���S�Td)"idQ��2.6�N���XU𵋅�$�. �/������	���R��� �3+� �m�ܶ�6Ғ��Gpݾv�7�spN���jVӌh���7$e	86����5��/���;.\ʑ��RD�bN46�Ҭ�$=5/�ڼ�,H���6�T��]?r?k���w�����	�qxz�z���L�D߱���*�z�jQ� �|���e��mA�t��GRb� 4K�����T#�N�j����Zr5�c�x���;|�*�����zitL��r�a�ܞ�x
/m-p䱁����s/��F��84�r�Oט���K���(�\�Y}Xk8z�@��h�t�t4��@�L��%��UZC�{v�p�{Z�1P������\%I<�j�4���;��]�l%��1��J$\�y'(���v���zNYE#�J�4e�� �� �o�����_|���(���0+�!�Xm�;Xߧ"��,��j<ʰ�E���W"2ǰD�/0Knq< �w��w'Խ���3����^B��vJ���kr ư�G��P���=��w�|YEn�.���J!��B�#�{<�b$r�x�^:s��4sH�*rH���0�/}�ˇ��!w��'��t��f���8m{У�ǆ�l5��42eN�W#�L��o+;Ri�8����e����=Q�roK�];���b�f�S
t�ۿ�5��O仟�z�$�;�x=Z�]K�4ީ �/Y@4!�k�X��w��{�Aqj��0�02a�#Vaq�*�Yyz\��>���u�co�[:(,��w����)�]R�łM �
�m
���p!�Z�aᾹ�t<G:�p��w�Aީ;���-�����E���ZOq=��N�KT fV��<{���W�fk|������6ˮ��֧�)U���^:f����#絞���2��ɔ�����lp��aN;�I���{�S%/ɕ��{ރ�#�?�ā�..�<j>B1�H�ٶQop��ypS���n/�am�6
TA��lv�ҭF��)M������#Z����h�D ��lde�}��6��q*�Vx-	:W��聍�9��n��:$SRgUy5��� �bx!ynF�(����W��^��㎣U�B
�v%t�	"bE$.��=��Q�����B/ֶ "�#������l���m��lG����o6�5-��33E��I�5fY]�dM<2ۯ��[�+K|��'���wf��}�ZF�ah�|���>�<�n�(���vߍK���J��<%i��;@u����x���mg#��%��]n͉V ��}s��h�2��n���p����%��r�f����%�f,�A�IT(%�B%Yz0HF����$��@d�	>�� �.���2�-����R���רHR�I�Ծ��r�]Q��&|��G��9�#mP����&-���H��E���kM�q�O�h��2����kBz+�	f�����U��5�0G3��^s^Y(h㢢u�6�y ��GMid�'
vY�|R<��I�qTTTZ�<��7ӹ�Cu�U���gbJ��A���
���F�(�k�gJ��vuF��;&}M�2#�g�ס�*��ݡ�]_�Ԭ�ܫ
��%�)h��p��F�n�y�9O�^��<x�{�[)Dࡍ{�Z��x��=G&q/'sh���9�E��T4�
Y�W�w�G|�Պ�|���9z��Ӣ>��)�b�w1�,V�6O���衿��K,������a�u�����3��#��� pc�!���X���_�G���4���]h%s%刺hD��
 �v)�ڙx�@/�K�/}v���2�{�x.�W�y�L�>K#�M�z������+�c5���+�"��k.��\�a`����S���L��C��y��]�����E�#BM:e�I���E�@��!����E|�0Yx�4"׃��=�~9w�E�����
W�(�A��8u1���a^� y������h r1���G��i=at���	��\�߶<=���V���� P��	87+O��jʨ���6I��_�v�9�0����0�~K��W�t}.V�C����נg�>60�FL��d~HA�3xD���0�Ǩ���Z��b�T®�k�R��: �df%�}P�a0c=]�@g�ʚ��)�G\��k�S�=WQ������Rs����Æ��&�\��3�0=��8̬�Á]!���� �z���g@h�ݶ�b�N�Eh����47��¸n�ui��o��G�P�fxٳ�V��)���1�gR'[By�a��2V\��J��P����\�Fc�̛�|���d#��+)oR�����͂ ֱ�zz_���`3�m�7�P�<�ѿ˞4u.�[�_�\�Ӌ��{���)|��*��&>��v'�~{@ځ`�&�7~Y�Q0�k�8�&�]�B}i�
�:�O�S44<f�p�u���r�{ s��ț�f]�ҩ��.��]@��7�唨�dR[SY�ǗF���@��(�'�e�?n���Mu��΁�� #��$;��U�xÈɥ�x��{�Ǻ���5ן�Yv�����Q��aO��@9���j�����\-�6bY��vO�]��௱ѡ���W(Oe�`��`r�-�|�$�Q�65�v���U�N��0��zY�S�5jך�s�0���o��%�oJ0��e���[�&x�'䗶��V.4E��:�P�2��@)|�[���ab٬9�C���8���t�t���Yq3��@Ȝ{�y�Iz�F�u��R� }�������� B'�c5��SV��9�,�BzX�Y�*�V�r~^�t��f�}0��E�~H�h���њ����O�_��s��+b�
��ݠ)�y����W���0Ҧ�ʢs��e�.E2�|�R7�C�T4n>9��S���a���<٠�r��k��I%��7Eר�!�5�63�^�������N��>�}s@�z_�Ȗ.���|�p�+>[�Z˒&��=�d�.��-v�blϩ�w�e��.ށ��[%B����\n:� ��?X��^fI#� !2mA��g�w|��X���-r 5��VӇ�[Լ�EbM�-	Ii��⧥tp�������I���q�G�g3��Mi��H�J5me|���O+\ٞH*��>bG��M=kϓq/��*�"�e��>T���`�"h]b�\��ndV0�уnY��@�u
���6��� ����H���l���d<L
u��`�+b�S�:��4��נ��k�4�(2�g��|-w��?|�n��Ē�[�jdX�����F\�$���'�-Z�u3tA�W�Hr�m�#ڹ*�ڢx,!LC���C8�i��4�D@(�g�la$�Ð��3H���	�ݡ���(�xt�?��K�����^J貇���C�/@�ӗ�C��C�Ka�Ć�Œ[avBjN>yP�$�F���ì�����+\��7P,б��	{%��O!{r�|�ی��i���a��쵗Tl��s���C^��]g�vAr���o� ���EQ}��G?ⷠ4`��\pQ��3��zZR���Q�͸kH盓y%@�x��F&�@��$hJ�*3��!�ɬI�XM��<�dqo��T��͕�OJ���gt@s/�Ӄg�X���eA�5SW�5�wƓ��O��ݽ.��G�,�N�&^�â}CYt}5!��Z�в�[p�)!��l�2@D����}
��۟����D�n���=�Doa�JO?�0N�&��1^�[�}+��B�~�����V2݆+UlTX�=�f]pl�`$���(��(�"-.Vn�I+�I�2I�g�^�;A����e�=³��^��r����i@p��h+O0/�К肓z��E�/��D�K�A��䥋�_q@�)LGA�5�������욶�ƹ�2�����>Cmf|��dpW��Ϋ��G&k���R����!(�#�������.�:������NS���xYK��G�*�M`k�Ց~4���v)���(�>��t�*G�|{�%�#�P������̻��u`�^�@\�sJ�4�s�1�CG��U���B�>���n�IG}��wz�>/�����"�4.Z�5�i�p�r�P�|D���$}��} s�"Iσ������L�<�	|T�Δa�5|kƔ��2��LL��%O���$2pC��s�k��b&h{[Jq�c1<�o�,u\�)AC�|s��=�x�I����v������[�~���~�>}��Z"7��@m+�J݁��0E:����J�g�|�Gy��z�d��/d���\[��ng�Y��Z3(��3�{8n�����I����[c�9#�ӯmsɓ�ō��<��?$�����*��J[��<x�(;VPx���񲥾�����1�"��'T���!s�m!Ʉ�}��u��;����8H  ���(^�NS�(sX��~o< ���H��=sh�l���f�%y�H~L��ڤ]Xs�h8R��@����<�������0�����-�������h�yE��V��j�b%.y�g��0>F��5��ğ�#�#�W�����ơ�ʳ\N2��~8?d�t�$���𵚷�2�X�o����;
��Q~�V�AZ6���p��������2�H��Ȉ�aJ1�ǽ�d��s���jG��I�?'���'(����a��0]������q����Ih����R���S�BO�$��[>ݖM�/���' 5x�l��g���"�d��~ƾb઼��@"�YC�8���q�iΙ�{a��?�?�03�"|��w~�Ӣ�H����G�5�5���D�Dzd�F**t#�]N��;8,Q�r�Ng�1al��ݜ��a�����B�=�E�?B��� ~��x׆�N1��MWr�w���t��p�+��G����׳�i�;�H����Ea���kO蚳��v穴�V��Li��k�K�Q;����.�@�qf�J-��xeh�o�
�+:HDD�1�>o!�R�<�#gd%��~0:Ķppa/�]�G0��8NQ������"�IY�xB��ۚt�Y����|X! F�]gK�C�/1k��/��]Ó �����.�~����>�QBq�30sp�mlx��G=��
J��2���*#L~ݽw�<eMMv8A���Bఄ����ڨ���bV�y��Γ����_�`�x�Z�̺��.G	�}&K1r{��C��4��g5 �Q�q�z�`R��E��C����U�D����������T0��h�9af�1�u4'ƚ\kV��xS��V󀉸�E�ƍ��HW(W��_
l������]+K�w�kyz	�,�lә��֒'z��c����<�аp67�t���b�It��Ġ9��r��bYB����;�lT�oXmS4:�ڻQ�+��oMy+���Y�0b����rP�T.
}�fh�.a�W�����v >7AYU;�����|�t�-%��@l�������j��^xN�
� ����t5,���̓�=d��ڞ,z!�l���R���
p�X��^A�or�#`[���P�<^���><?k�C�LhX���b{�]�������'�a.K̀^f���j0"d�Z���?ш��,�/�W׬%�V7�"����%F��{������BX�� F��Ϳ9�.�C&�f�A�ӑ�C���E�Z�������R+?)�Z�5�q5��¥��.��M�,�'�.%��)�[:M��K�G4��s���3��a�S|p�5wS���[�x��1Be�ӆ{�FQk����rm;(ب�H2Y!/��K�u�h�c�T��i�o�݀2p����	/����B��0�����Cx�p!�K�Z�3pw��n�j)�	�������3�ٍ�*���$�6�7o�o�t�������;�L��s��A�J_�z�n"󌅏��s�pXq:a �M����+ڭЗ� ��Y�U�t�ħ�>��=Pι6�}H�o
�{0����z�Q�F-Yr�TT�	,��:���$���}�����Z��d?
%Ml�NFS���v��1�4���L6��%k�f1��5=��>7���� ��`p�t��R�ZR��ݴ�Vpad ��_ÕX���aO�,؃v*��+��/=5���ݧ��ß����s���Fɺ��$ʝ���;�G	/p��Qم�G�Aw��,ȑH|@s�D)�ޛ;萱��S�.H�͖N��+���������W�����r�n4���÷������d�p֌�d�N|�/; 5�z5w�
t���p^�5>�S�9T���^�2 L�{-�Lߠ�Q�}|u>/�n?�ʙA�	�ZN`����;�@.�z-6�|i7��5# A���a)�_�'�3���$!S�]AB�RC���0Uޯ_�"����Y~Dp'KeEX �0��D\��c�t��؍��AY�Q���`Z� ��3�n�`,U :�O�@suY�Wo)W�6�>u��װ�C]07$+ s�H�D�G�{�����n.t���OH']V�kg�*�Kdƪ�K������2���	��M[�tb��[��)xƂAS�q�|�z��_�����Z۾�3�(�i��͚�`��P��,h��!�v�;7<��s@i|����W�v�A��	>�O.�W>E��I�����<�H���I	�Y|ll�>�6ur����>?��`q�U���k�/�[�ҭ�!�.2"E�-u�Q�4)��}F8	��6UJ}�D.��Ǯ6��H�l�H�
N~"��9r�m��P'b,�t�!��<�kg�CA���l��迅���ew�|����}��E}7���ٺ��a���{�xZ�����o�D�Un
!�Ud��&gI ��G��-���4 �_s�T�>Yw���X�W�/��U5,>=���[f��d�����aY�f��-�����X9>�M�<�f5O�n��?�R������'?�+�3r)���a6i�"2L�)����0��Bd#Τ�u�f���h�w�Jy�9������lw����C
�`&GW�CÃK|
����B�K����n\�%�,�>/Ԗ_�@EB�?|���P+*�bi{�+�2��p2�б]�I���%:�9#`L��0�T*�&�ЄE%Y�`�E��~{yL�<jXӚd�_�4���v�2�ʨ�
z��]�K<� D+Ĉ��� ,��aA�M/�GzI��U�Aa�l���=�!g;%t�[u�T�rΟ(��-��n�x/��Y��J,�^�J�� �!��J�.�1H�T�|�(�]��������?����lq�k|%�h���<��.��Zg��ڈ�}��]���������twmI�j��� ���M��(E���-�ND��(������R��
��Q F<C֌3B�/��C
�4ɧ?��`����މ�D� �3a���)�io��YVI֜��>RMhd�YH''��U�	�3�r���C���A�H��ɗ��-���l#���a��	�Ѳ�8M�Y�>��k�͵��j�ۭfM�x
v�Ct�]�CZbj�Y2��L����3}�2�":d�����_��0z�eH���� 	�e�lD��ts+,q"�'&�a���Su�d���}��}�-������.���&�Ji�`W��1J-��?C���4��?��/�c癴�PN�!�2��{z�UT� ��8��b�p�W�򘝕,��!��4�Upc�àD#)#|6;�@ԍ�I��0x��D�)D�`�Bu[C|Òx�z����C�[M�O�%�xS%xyh�0���`fx��&N�f��JhE9�a�l>	�2
"%�:����|�\%�m,F�l���5�'�{�r��Ƕ,/FS�jE���v����+�����N�������3����s^?{9�dIKf���X����Г��S�SD������a&�?[�D#���=檧F �NB����0^x��]��\�n{���38����J����f��U?͜g)��K���$ .:�Oúk���D����20�b�_�?�Hd��uWTi���L�/O+��O�I���佉o�"�r,�>�uF�~	���M\)��M�[� '\��
� )Fm��p~n���
��f�&�q.�)�ı�c�\�[j�)\���*���k�J��MT�Eͫ��'d������}�
�Ҿf���0�F�_�<�yx�3��k�ų�H�+���ӧ��l��Ѫ��X�=�=?���N����s1l� ��;�f_,��d���A�Q5�}�����٪��H6��#�����#����`(�wP�9�n������61/ -�T�ɮ��v��!�����5d*��o� �D�K�}M��tW�~�@�W�Y��B��� ��C0����as�1xl7���P��Z&�w
dS�-�_����x��;��u���K�+���3E3�GpX���_��In٧�"�H�딎��i.��?��&�����h� '�E��htpl�/w��U�P��KzD&h򚭎�F�Z����������g�|@� ~.�!( ���b�	H�&���#8{�x[ح���s���}I$o|@N���zc.B�P�>u��Q��V�I<�5��]�8�|�mE����VM�]�����q�-6���pf��54{�k��oy#ʌ���`���2i���/����(g�����{t�m����my��u��z�G���%_��c��%��s�<�É�Y�`�~��������M��M��if(����q�d�"�'���F{a䰐�ƒ���R\C��=�Gmm	�!����?�Tk�G�mb����b��Qmg�ޟ�m�:$�����ƚ��Gj��b�ז��!����j�8ڼc�[�"\���o����H2����9�c��[�w��b�_X��bCW��#Zz�	���$ꫭA���QJ���{a1h���.�H"�����!��R�d ���O���j&��6"BdQKG��h�V���ry|�d2}l��k�,�]x_����a�)�yR�DE�D�ܡ�8�*�ď����HT�#M.o����iE�{�\5������<m
�b�,K90�	IH+t�켖[��`�黧����l���iܗ�AcJ��[5�X��0yc�j,�#���$����� 5ɰ�7;F�6�Φ*l��[��9�ݏ�߯�l���Y�W?����|e�9�R�&n�I�w_A��g̢kՀ�9抚���: ����7��yͅW�x��=3��;n����g��>[t�i�OŇr��Y��%���{��M��ʻ��ǭ���;�Ka-��${@�]8��\�2��6��zt�Vch�҂�����z�yyK�Y��}���4�#Ƅ�v2
Ι�|��Z�����p�2�簨}��ǂ��Ka�E�d�~q����K���sN��S���l��C��.�x0o�s����Vdu�1������&IO/Zh���`n*E��x]��ےϲLsx���
�v�'�xa���Z�����o���������Ϧ̨y�w����	Ĭ��a��ӛ�{����B6����;�~��gI#�Y�J�]�W,,:"��voo7��Z�VI(��J��-�D!�b���1��O'�h/�sm�l�*DM��?��&����2LĘ��㸋p ����60�m����^�)B�ǉdY�}�ԯA�|�n�*O�6Y�Ȭ)Eǌ� xd������s��aR�kY/��pT1��A�ӓ��,�z�����z^�W/mBF>�2t"�����]T1;	'gqw]r��b��k̢��)s�?�Y�K��|J�z/~OD{��}����࣪�'/Z�|+µ��k�K����y宰�M9�� ���n��^��H�Un��C5 �W^u�,����d+�i�PS��&�k�Px��ˁ�Z�,�k�A;B�;WL&k�+�`��/qi������<�����ި�#��G�H��ɟ�ʗ�ޢ����#�F��HX#J��X��Wt�c:Ԋ��(�Q��X�Z�EA�l��FTco8`�:�}L�a�յ7�γ�4�".��p�V����� ������֨C��UJV�n��'��V�}�O:e��z�J�iF4k:����P/�8���4%wP�a���W��[�H��r�C��H�9]ŋ�EA��vG|c��J��v²�`��&�"����~ai����쯨G�f�L�v�So٣��64Mu!�HeMȄ�ԟ���W�ٖͥ#�|4Sp�U|�(��e��{~��?��;�I.��pXFפ�"i�6a����0�!;�=�($��P~',.�#��4���k��1�:��(Ҳ�z���ӿ��ꔩ��M��j�ﶹ�C�*RݶH�{rLV%�I��V�͙>��*��o�'Tx�Mʩ��VmA�)�����a70�d��<!4�������+�P������JLl��DY �\��K?�u��VFl������3�Y������c����{��	ǳti�vi�5��z�/j
�v���~5R6�πE'��̝!�q��!�׸g'�|���
�ZNb��#�ve8����a�/hB�� �1�n듋���
F���x��IP��Fy@ɮhmKX���[v¾���O��8Z(����A�U��Q��~�I<�yW�ڱ $%}>�!>u�o��!(5��6���z��,hu(P��=�6�`RA_����g�ˀn_q��j.��q!υ|�EpT�,�[�^]������É�(%��P���_}��FgǙɟmFI>a*U�Syh�]������>�� ��˵d(�5+���cEG���y���D'�SC�@#J��z?ۑ�I�g�!s7	~���"�H���Q!�R��n��$�pΟ9K<)ҋ���y [�$���wϿq�<
e�z0�<Xjq����/γ���@�y��a���W��m��]4+^\W�����7�\z����?�KY!�Pnي!G�gzH^���#d�S KG4��<U�,POցv�o!Jj�VA�"�D��W��-�՜y�]��x��������Ј��$�ND� V��fIE �ϧ��&����Vʳ뜜�9�T�7�+>׺��H����c/+p�Si�\)�ʦ������M2F��ϻ+AR6�G!��+�T���}���?byjwM�ɪ�[�=
&�^���)HBi�
6����YC$���L�����<l��l��5�C�ܪ&ڽ��3"9iiQ��,fO����C��ɺ4���I�y���g�T3�����:��m������	}����fMpe2G��8r���:S�q[���%�85�����9�3��m�ο:Ig�KŤ4�f+8Yp�@u� �E�����9%z�������u�eU���	�c��jM�� �=2��,ok?s�,��������K�a�3ws� ���㓏�%s���%1`�m�n�=��"���X@ k�!O��쏙�\!����n)�DA:��;�>,�����I8�)J97��^�U�V6��k��kVgN*Ff���x:?4��Н�&	�eO�#���Ί��`�����$�p�m��Avtw�y`�PX1��^Qy�,װ�6e���G+�Ӈb�'�ґ�X�J�,��3V9'����0���Fi�%EP�d���*�7B��P�����c��@��Z=e=��O�<�#ǀb5�r�#�Rܘm *��ି:��f@�Jp�l��e�W�ҬCv7r�kܐ��$"�k�:M� ���;�r��"�x��A�#@PkՈ�.䦹����{��T�PŁH�U[g��+@�@��zƦ{������J+TC����e��� �N��k���0�ɠ��5?$N5(�u\�f�f!j4��q��'�w�v�M1o>��W����Q���	-�I�PVY.1Udk0�K��ͨ�_ǐ~�M���1����j�A���cs�`t�(�H���Y��)D�{̺�QY�-�o� ߽��t�
��!����` {_U�X��<���CM����w��#^lj�7%���lK���fS&��c�4��b�]!>=��0~�5bK�ɖ3#�S�d���[�D���'�(���i)U���x�^.m@�?��j���>:w2Ͱ��IY�Fl�)8�(N��ӎ�
aI��wX���Y'>꘳?3�}����Z3i���E=�?3�FÐG���~�j�Ҽ��!q�K!�>����o��D;��P��+y'(����B�L壜r��OFn�s��|�jZ�tĖo3�
r�?b��Lň�6œ�j~��궫CG^��}6X:�d۳��u�Z��rǮ�q�)m�;��$΄J��K�*B����C��F?` ����,| x�fƞBl2��24�YQ,PR�Dc��/ �=T���p�mr�5�?�v����U՗{�{�u�;��g�v�գ�@��Gzuf�I�ywGs����:T/�d5W2F���h	hp:d��)�srzQ�ׂ�'�P��.y|pXY������6�����tεF�N��V���L��:�(�w��G�����zu��t����2�
8�~_��U��>ج�U{7C��J�$��vB(ls���a!���`��]�5~)��pP�T���PϸK�^��ۋ#���)ߗ��1g��;�T:X��PA�G���j������N�\;����Q��Ȱ���a`�����6�9���=L��Ӎ�i��F_��Iw+��\�=����qJ�iH��1 F
����Z	��n"-�HY�K\��w�@O{X��� F��S�fp�֥U��Q�����V`��n6�����'>Qg������q�/X}��[EH�"�U��v฀���+91M�f����ڇ�$s]�3���9`�X`��n��E�T�iK~���(�?����d����
�S�m��VM-����$�Y[�F���+jK�*b�q�^��J���2{,�54M(�X�.��{軰����G[���#<��x@o0Ϭ�g��g��'غ��ngB�.�;\���o$q�����g�z#W5�������k �}uWߛV<)/���ޤlQA��"K�AA���@�(��5���ˬLU��v�A���$G�k(O�+��jA�� ��\4vw����ԏ~�X��} k�9�d�?'XWL�z_�
�Y�WwH��5a���8d@n���QJ˯���[Ԛ��������'9k��j�xHN�m�%�'^%h4FK�G����đ�gw�jgP��]#n2BE(p������[l(�*x.�nw�!�Ui:<V����#=��ޙ>�Rvh��'��w*1� ��>�FKd%9�$<�x�X%���ϸ{��/
.턯�/uY��v$���{?�іa	��}ה����A"_��&�v|X� �e�D䫼%e}�������[���$��̒u���:�����?���G��L��A��XWVH\��,�-�i�>t�����vWp9;{�ύ��c�'����J��]�8����Vi�.)ĪLAX���/q�q]�2>N�����}����+y�9;�Ō�~mו�����h�a�y�t0X����z����x�w�&���ukʛU��Mˉ����V�6�%�}�6�Q58��~��!>�p!\�������qy07������l]�)���0ۺOЇ��NOdo��$>07o�9�I��6�ikߘ{O-�D�|+H)�O�:�+>!���b��D��BN�&�O�d��	�q�c��,��\��<Ul��z��a2H��"�C���Ug�Jt����}i��يRvχg�=�^
�2M��]�k~���2L�l� ��A�g��t�{4���qx�������v��>��b���J�`dR�̛J�va����-@�m[hH\��c��E�I����+܊N���IH'��k��nr1~qA�D\�I�b�j�j��dE�i0N�F��|������� ��wt��Vg�Wg=���w:�~��NkPc*C��
;�|x���V
pA&,#L�>V����Yp�;ea]2�,V�IE�)�,���;���!s��>4��ee��u$��8��G-�3y��g�S�ш٩��Z��J���)��y���!��Vt��U3Δ��APz�^~c��|�L=�g%�]���Rhg<��ORIs׹ǏB�@Z1��N_�b
��2/��F4�p�{��/A�uV0J7���k&Fc�����f	�drQ?�6&gT�,Ͻ���Ñy}Q�䒇W��Gč���b+�z3�&Nȱ/���4H*���O�b�����?��Y�~����/\L���T���|c�cC��H6C;M�����8`��X�o�bՃsn�&�C�W�SY�O��z��g��b���aɣT�@�#���}���>��}Y	��#�|OSA;|��~�-[�VԖ)@(����5j`sk�n�E(�S֭2�Bƥ�C�������ּ�d�r(����A��A?�ұd��Ҧ\l��~�*�yTf��[jW���]~�{0a۩���PG�GiF9���hC2�����r��_�����`�L*Ё�H����mfy%�x��^����M�g~9{���Z����<c*.Y�[�I���U�T6���zɏP�z5u����d��}���s����⏠ �W5$aa� �l����0jv���F��\V� Y�2��2v��3��*ƃ�
��]F��.%w������r�F4�x��<RErV��,I���Y�Y��n�,�g��(\6oUb`��SkH.q�7�n+RZ���z�� P�ӯ��&1�~���/�N����J#ez���d�s�s<���(�4�!bw�)7izp|�*%�:X�������s�b�p��:q�򈢵V����!q~��S�к��s^�5yj����H�����wPt�q��U>H�H.��=��P��A#|an����=�E���deL����?����������#�4mi��g�M���J��bW�����G6z�`#|�[��'DDg5�(%��ZMW��� ���"_�_RR0$�b��r_�7���� ��V��h-s~�Y���,��;Π��O�n�$�0b48Y.�,���@�Uǈd�v����\|`Wo �z�G6�l$�Ʈ-�v�,���|A
E�9O��]�2�y5�+���(��^��7����6��h�����OZQM_m��/5~2�]�T/���Y��:O鴹_K�C3g'�z
�v��7�@�Z{Bp���&+�Ő��M��O�}n/�ڢ���Es��r2l|����=Bna6y$$��꽛�^��Y5#I�� 5��f��a�X��,ddP��BƍՕs� ws'5vC�Ǒ�.ľt���["Dy2���U�K�U��8���$�PN��μ�Ni+q��a׆���t��/%{��e��g�����D��8���o#��a9@��;٧gir�����"�1�U��pY��T�@W�Pf�;�U�j ��!�~�}J7��!�����>c6�*�-�W���n)g������B�1GY���A#�Ўݙ%��u �� ����S(�_����a@ҌY4u^��Xɸm�ݎ1�ggc|^��qb�J����q~݌oO�yG��":������m�hd2�;M�ɣ�A��h+�iX�J/r�q��V��@�%ur����~x���_/���8�����ó-*�T�a�[�l���ԑ��ⱘ���"l��4y��̏L�%�e�%P�iO�>��Cž���ݔ@D����i��0�;��B�0�v�!_khP���6<��[�-He߇fj^��˓�B0�h�_���\_�&�&�k�f�;�gr���ْ���_[i�z���!G%�����v4��@±b�n�n������I;���3?��N$@�!d�j��F[�$�r�����zGd�w:�$��0��ô�M�%����AV�7UT�D�CU/%D�-��JZ�`K�S0���y��������Z�H��]CB������Z ����ujw0��uc���\2e��N�NQ��U��6|HC0b�SDn=|�9Yc8bmY�Ԯ�B=����H|i}��f�E�n�-���?����˅��2�A)7�겄?�d�ޏ�f���qab;�m�3�[��B;Ք�7C�&��G��O/��5H��f#��1ґ`(XV(��08-ݺ�ln�.d���GQ'�lB�J�"�ˁB�m��6Q�˰��A_K6�YO`�/̐���ٛ����#��c3��Oi̳�����)��xE�c�CoW����;I���T�ϪP7L\��RA����jy))mi2=�*��^�R��$��6G���T��3�㼅|�Q��/��v�������'�V��-�kKQ	��c}�[%�-j<�$�H���\1�VqlY��"6
�tP0ڿO��Q@n������a�Z��f�w����C���!I\�%��^o;������fcJ�Q�^]Tu��K4|x�^
VU���Ʀ����d�����g����|����d�a���,sy���h�A���'��F�~1;��
d֌]�)��p5�
k���(��R�r:+�
9�P���nŪO�BU�d���ذ��_����#{p����5 ����g�}DP*����c���P,���ۿ���g�:�پ�O�A3�]�kPX�Z\�F1Z�ů~6�<��"�7�~��0��[6�������G�T��}���y��99��G�֦�9Jc��'Tﰱ��}��U7m�����(�2�W��_C��_�����=�1��]��"b�@�"B�4~W��7��!5s�b��>�j
O����h�'�u�v�)��CX-A6#�&��v��lJ�)�B��-L((o��$�-Z.������<��Xe��Q�!��z�$�y��-^���m�]Z�PS:��X�1�W�6*�+ �Ɨ�����%��X�lJ1e�Af������5��8��UE?��#�Rph�R�t��x���0�p�D�E�A�X���G�������;� �;z�d���iI�?�_렷����E����������-�� UIzɫ��h �ݫ���ϑ����b3�������.d3���#�W������,�^R����f��Aj�#�=�@�`��L�C��3�뜻+nJ1�ֳ-�7	F�*~g��]�2~�dF�z�"x�Q%5Vc^��;�I�K�N���Б0�w���Vah�Ҝ/+�,AE����l�N��������-�6��	?��HO[�`Y�(?�ě�6}<�MOB��������"�g����G�d5���Σf;������Dդ�|�Ɓ�u\��?�3$�8��"-��s�n0S��m�w����i�nٞ��X��1�����Ȩܕ@I����?��u&6��,��f������H!N�#��@���Sã�_�
T��g�I���j�Qm�˹�g�V|Tl��H��Yh
�O�|���O�a�r$Zٻ�H9e@k&�R>E(.W�ޣ�~�2��t<@~�9���pr���UQ���Pg��DW�s��΋ߧ|�@p�?�bC[�G}uYo��7b�e�g ��@��v6�J|�m�}Qc�aK҃}��i�Ѩ9F,�p!��{v&`��)���v�!U�+؞��O�D$�5v�c�b1������HtKPQ������C�Sy>#��O���� "q5	�$^+*Y*nLLYK��M��,6�� �[A����6���.M��$�Ӑ��C�u�����(�
K�#�R�,f�l~#��lhO�����#�k�㻗�;�C^����0��f�KX�F�lC�X��E��\eC-g4SI�?q��Y���M{a�	���}�y�S��� ���A�v'~�ޭ��D�W��&����\�iV#�l���#�6�0�v�+�]U��c�
;4*u�ӳ}iY�,�)�)��
j��=8y��nRkgK0�����̷�Tw�4M�-B���i,^�)�"�s�Y$Ey�<�=�?n�ˤ̲�M�۶M
:�̀?v�mV��`=�	Nk_?&O���HEQ[�H�5z�`i�V���X��;4pzl��:GE��F��g�ļ��<����ڈӍƊ
�#܃���]�,r���&�^��;y	5��f�bKb��p��i�<��WE��Ƶa����$�ͿE����eݚ��2y+\��e�n�Ux�ދ��"��BL$J�T��}X"KCET)C��ҵg4tp��^tQ� ,���w�>���3�,����`sĀGl�7aa/�y,��K#�CF�?.خ�"�+f�8�kS!oCQ�&�Ўu+9b0�Ԩ�܄N����/11T�ߵ���<BU�O��8�#��\� ,�� >̾~Zq=(+\���w����^96�]A���4�H�}н�B~��ͰLس�U�%%bh����r�"�g>���q�Σ| ��Zfg�D�`�_�6�fPr{�u�����j�V8��Tθ+��m*m���=n�*���)�lF��?L
k�B!r��
�W�-��-�K�31ISb��� q���cy{�_��[�l��g6cE��ݖ@�������)������u� ��q���������m}hRxB�˩�a����7I2YA�و�/J�2⤊�Id�5�r�)k�%Fl�7s58�fp�:Ul�Қ��YTZ�Iq?���2�Q��?Wrkf;:��t������qE�,1��~���먘d0vR���\�
	��d?������scn����EP� �����J.$��L������e��;��O:���ȫu�:����L��Y���k�p�:!�(�c�p�{х)�}���kF���`��R���o��ta6~�L҄C��E�>T�o�6�"��RE���3^�+�&|��v$�����;r{�%pco~|�Y�'ȩ��ʭ��H��F��U�8��`!�kү��.�|���0<Ƒ�x�^��[���.��y�����w)P��5��SU����`��3֬$�1Z��]�*�t���цO�- cC�5�]2F�g0�-=m��6"��-EM��8�UU��󼶶>��T�e�;��>Y�K7ϋq�I�T^��Q^"GF�_0N���á�g�7���+�`6]؇��u��V��E`r�T�`�iX���u�Z�Hat/���7b��mc>�&*J�eйo`����ކ��蝓3	���j�W(4�s�l�3#Rw���m=�a":ߜɉ*]�~9�o�A�Hv/J�6�QDՠ��EL!�1����FpJW���G��YI�� Tb�A�ȭw�����*���F+Q�sA1y��<�����6�<��9�~9$-�z!��f� � ���❺��4�����g��v|㽬�Z��;(S�0]����������hq��&i�o�2#�}����4v:�[϶[�uHDB۽�TS�k�G�hCb��#�m�F#a[���l�əA������8gJ��,pO���0%h7��H
�ۂ�ÚB�Z�å2�����
c"��b����3K�@�X����j�9mc�8�;gF�:�y�v���5�َX��_��r�\I�ݶvQ`)W����e��7͌���N΀_�1r��=pME\�5	:�y���Ic)s%�^X��-	G�u/�5p�A��u]�	I�:����R����d�mp�c{c��J;�M���NM��7�M#�'��r�Uջ�SX���o�ҩ�\#9p"RD���@P��]4�m��C��G���3LD���z�9�e����Ն[�)	���A��YZa|?c:���v�X�������;<Za<�ԏ���*k���(EP6 ���@$�<�#�c�k�����U$�����g5ú��5J�OK���yR4�=���F���_7W�_GU�S��0��2��.Uܼ퇄����C>g{��g�r� (�R�L2-U�0uH�O�UW���=z;���v�I��0���b��8�ߋ߆����sJ�@ŉ�<	EQ�~	A%w����0�͢���Z9RSR�,3j��m���Th�zk���&�_�f��t�Q@vp2P��y� N�f����z�
0��
�5Aw�K�@��9��b����:�3ar�"P�kL�$!8dDT�u�/��Q�3	�+��Ta
�o�j�BF�ۅt^n�D�\2�hu#�V�{���}��H�9$�֤��M)��i���)+�V��b�U6�ŭ�{�lzϝL��<���X�k���C���$f��(2�������1#���8\t2�X-�ʊF�PR�c�p�N��2��|ȼ��B*q�]��;����T"��Mأ�̏�+Q�L���r@n���~�5MIO�n(%.�:g's��2Mn=��2����2	�5_!.K��]�ʹ��~���~��rQ�Q���F��_N��k�*e �O�WC��Œ%�1-k��j�9�i��R���$0K�8�����Z�j��:��j���Ćr��bt!\�>ǭ@)-�MA��b�Hșuw2�^m:�Z}gܦG����}EK����4��yx���F�&��T�����R�"u¯�w � �
e����wVV��y�m��{ Y:���1�gi�K�?���}"�>��H�&��������Y�N;�H��("�M�����lwy���udLW�L��h��M�EqF�Ӓku(��?]�x
S�`}9�������f�A��J����D[2W�(�w�>���T�鏛�q���ЊT�
������b�dMg��3L�nb&9��T~K��csO�߷������\�4�-�c�ɼ��@ڿ��2�rY����o{6;C���w�1�/�In��jk��z�ě���,��P��t��D)oր�f��g����W�������8t�eUI;KH�{��O�LtLe�*	��gyo�{������ �T m��6�(��s��ٛ��S#��&�Vf\�2�{�Ԑz@@�b�C���)$���&�na�[�!�nV�����ae3�f6E!ɕ�mI�H�ln���9���#�����0^tU�2n\*��|:4�����^��c��YY|���C�q����ߨ�T~޹%�����xx���/������5�����l#u=x�R_��ћ��-G��i՘�<�0rvZ;�RN�$�u���� ����3�]�+)�Pt����2�/ζ �
O��5C�Zխ�ƌ{v�A�B������{��V>w!q�V�ݷBf�8�;�6h<��{p�W#m(�@��*�4��ۏlW��(��!�m��h��AM�aL��VU�)��fն��8��dZ���ŷ sL0Y3���s]�1x����Q��O�Vjˎ��!/��:���{ӷ�� '�h�K�e�?�p3h���q�V�~�(�d�j���O&�E�+��:O�����8m'���	/��g��`?�`k\E� ϱE��e~�T䴮���w������xZ�x�? �f��X�m�����ptz�\�߽u6-v��w��kDEb������?�[$�xܡ̜����ď4�3�u�8���
5��j�n*
��:"���!�:*��qO�C�C^�Si#�;���@E�D��ҿ�
!(�8��ᇚH�[�7{�)��p�|b$�H�
'��H�'xv i��7I��R�Q���9kJ.}Z?<��C�>�8UB��2�n��;h_��=�t�Y~���\hSm�̻�Qo�_��`~�R&x���H���&Z�KD�?[ܬ�+�<�
�˵�� �FF�n��zV�E���ˀ�]��<0��Oi���oq��$9QyXź0�$��/�d�1Eˬ�e�bc�v�痕�Ђ�Y3��Yu7|�ĝ�0��)=/���!xq
{/�������+Ǹ[èS>o������8��,������b�23ՠ�?(��Ӳ\�1w5�_�Tla��.�
Qǿ�
@
g�n�3K �����n���n섫A�[[����@�
=���o�)g4��5��W����y[e$dXH�����5�W�k|���.x<	�b��@U�MŔ�"ճ�� ٬�W��(�E9}�����p�Zq\�&�WPv�^RKQ�j�)l��p������p��� �� ��jG�\l\P��&� ���}z��sܚ"��%%�Q����8_��;D��<ن8޼�Y��X�h�֙��7o[�
C�{���]� ���pA��]�]�* wjMP ��N��m�a�Z��ڂj�i���҉�p�����-��l�Y��l��6ɖ���H>��D��2��L�-E֗���u�5�	�G�ri܉�M��]������Ί\Q�B�����^6���ȱ��)]�B�>bX'��n�wG�������c	�٬���n�Y�h>[��J_?n{+S�����1��3�.Fλ�����$Dfb��n<��YC�,��~
�`$@�{�TA�r*���xI��F��	��B��Nw;Y���]��A�|cL$�UsH1�T�R!�?j�.�k1�8	ʽz�;Fh�z���:xp��
}R�z�l����oό��7�$�1_�W�EB\@��7>je�(�1��\��뛘��{V�HՇ$�j�͖��*�%}��nRp����q�#�mØ����z��f}
�~�c��
V�K��l��P>�5���p�"0Ìo�(�L�K+�J< ��SD�]*w�C�n�uYT����x�4���Ck��U�ׄ-�f�� ��;QHa|�C����Lsk����� =��RG������Y@ V�,DA�F�ٲF����Hj����A��;7\��,]T �p0rli����}cS�tE� \=�+h_}Q��+�ļz��p�n[�&���;kD�_�������:"�=?}�+�f�^�j
q�������3 ^���g-�	��m��m�����KCZpW$#���3��9�Vm�n �Q"5�!�3����lX�c(7��A��t4e)���^WM{�B`[�~�}�sOZ�$uO����rC�4Iw�Q�)�Q�SW�d`�|��"��4���\?E���VI�Z)eUQ ��\���1�-�ѴQ��h����F�����9�Ȯi(�vK�P�ŏ�%N7d���ޑ�F&���^��W��߾�d߅���M1S�e���+='<u2�-�{H�jL{���$���!�6����6�����Ϩ �� ��,����>�d8y�84Y�0��/���;*HcA+\+���0��_3عF�v�����)Y�A�$�Cjf0�g�Mh�%�E��bR�aXb���L��qa��c�y�\!+5{�֏��]�*�W�gH_���{b�ȐVi?EJBZk��r͈ct�wv���ż�>��0�с�м�ޙ[�uj��u3��ǳ4�����h�ܶRɎw]$x6+"bЪFFS�p+e�'��kr�r���8r=e"h˨VU�օCh�4"�[W���՘5\$�QgC�$&���{��m�NHWp�H����FXﬓ-r�N=�V�����*uh��!��$����F1'5 9}m���W��{���0�C��b��	|H�׳v��d�1P��Y��Yy��P8�Uh%Nu� �� KT� ��+��!Δ�R$���7r{��z]����"�� v_m���� ���7Ŕ�.w���|����'�ې�=�`�S�|V���������{�Q�R�CQ�B�&�b\Gښ�M|/>�_��6������*�IM���{�� ����b�����/~�f�xd1u�F��<�f~:�Y(T��g���עz��w,���@p/[#���*��|c�0 �6��^�3ՙ6)_�=q4���5���~t�c0���7Z��k�{77���n�p"�{.�&Ԇ@[�b[DD�x�M��C~�z��M�)��fn]Q��Fxtr�V3���|d�#6 !�!h��E�僱i�����O����%�MA�Ə|P8ښo����%�2�k��D0��5y�|�K�7*Kѽ�-����ԟ��&[�yz���M�0�e*��ow�A�����B̳���S� �a��3��R��S��������!$���M���坛Np����_���/�NGy�}�z��o� ����xdDO�@j׸q1�'�Y�����p
�+����3�0:��W�:���+��4�4BQ�d�"�o����/�?U2.턅8��QR��
)&N�e�q���"��lnl�\���ȅ�����8�Ѳם@��Ja��G�:��8-�G�>�
k�g�*�B��L���"����w>й[c�؆�����;�V��OI�%�O�A����c���e�{.W^�bgY�\?���������-�Yw�(������7F�9�wq�1jw�B��,��r��P�I-�����J�u���%��8'(ff�4^ � ���@�B�GƧR(�����2@�X���3��e���A��|X8�ݟ=y`��}ߩR��b��?���e�K#Kk��F�H�^�t�͓��Cb.�Q�T�؅��X��ľ�_�1��GŸ�,N��O��ޟ��[^��
9��/�;��e	d_�p��آ\b.�9[kܖ��d���$1��'_��d"R���<�]iҝ^JC!sn������6���K�l"�uۗ�"��٤:�-��ۚ��1Q��Vk�Q�=���5@��aT?VO=Lx�R�@g����7
�� �,��=�b_�S�%~��p�n�����|)a6��V�������i��	g�"���J���v��F5���v��J]a��lp|�'�V�Ð��ɮ��?x)e;�_��*26����p�`ZN������j��m��W���@���1�R	�9���3t�c�N�3�S��*���z�N��Iڔ�<q�h��Tн�����́�Կma���xÎ��<6����|.��DU0�Y�l�bjo)*��hYMP��W�q��#`��~��2D3���< � I}@�+�Dn����9�%Tb��,E����[ṵ&S�ݟ��f�}����ґzXحI���D#��1r�j�te9
�k!@����)�R�����k)PT�d����.(*��+�)�0�$�}�J;_Gi��)]�;LE��9$��W���Hb
h�(0�p�>�+e�H���ȮՈ9V�ܡS��Ӄ�	�3:��f��3^y̤����P��k��:����$ �:${�d;��a�#���s??2Յ�+Ic �3�TT�m���5�&�Q�e,��ܞ$��+=�#̒[�?����Va���{e��f	�ٗ�M\Gj�x�<8>�p���ҩ�*Z>f��n}���E�:�r���+�����:��e��	���a��tZVx�s��,N�+6�O'���Y�9K�q�@�>k(gӳ;��c��3�uL��v��ZB��o�g:;x<�b8	�ͷ�n�� ������XT*��"䔻���lj*:�.���75���+�A����S9�tW�T�R���M8@0�J:mNM�q�+5��,B���y�s�\U�11��H�#g�nW\��F�w�����;j��S.j�{��Ǹ�/E	�DAX�̛؄�'/+�Kx�'���U?�� RI��yla�g���2+�!���پ��E��~K�4�U]G�h���!����R���s�ʹ�7H¼�k���WF�J��ˋ2�; ��6��v%�y��*%%����j2�B�����
a���ͼ�낸�A� ������zBy�s�l�+�jDk�@3�_����
��@蓨�^ܟ�?<�.4t�e��K��{|��˟������ׄꗴ�j2pZ�=Z�c�X��f�>U[)� E��:�kd�k�#i+�QK�Q�V7��~z����£F�ow�K]A�z��Ys3�����떂	K��֧�M��͔�n��^Aх�RQ��f�ص�+���T�������7!�qҧÞ̆9Y,E?��4'��!;��b��ʰ��Z���;`�Ϭ�=�YG������:͋-����c�7�ud���q�Q�0�u���(#	�0�]c$
�[#f�G'3S9�5�e����Y�{�Xr�]�1Gwn�#t�.T�24�CR�kI(��h�që�w�OKL�6⏬�Q�z_ͩ6*�1'���G��8�Ҥ��`��/��[U����*$&Y���4㍡����"��B0���UAc�8g����YJ��v�0����K����]m�o��H��TjJ�Ŝd��5ݷ�״� �6�daٱ�d�!g�yU�j���Y��g����f�V	ѿz(֘�h���5��P���U�K���\���h��BdЁ�!h�.��T*Ώ�_��tq�0wѕ�H��i��K|��3-��壸��TQ��`�yl�O�m 빃�[�;�~$�㍊~�>ŮJ5f��\�r�G�@�{+�i��0h�F�0���峅��G-[���h�H����9�`8E�n*�!����Ƕ�w��w>���	n�����'m<���$:����RBsm�������?�H|��Jq?U���R\W$�/�4k�@	��ѿ.��z��l�9hkŹA���ٯ��lk��ˈ~�A[��=��t� �9e=�B��o�W/Q,����X�n���������Sz�r=� ��%�`�w�舚t�y���f�\8�Dj�0g5T$cL95�Rr߆�,����9N,L@�blZ)�'�V��▬��q�ߣ3U����K4(F9r��4ץ�
Y��	����)l�S]��VSU��"��{sP��M&\��S;h����vME��SF��8�N���H��J���"�%p�����Q�;��������"��ɓ�O�����@��l�_��ܧz��^%b?Q���6�.N2yǐ����>�Am�t�=DP��o�-��ʶ���RMtO�(����NP5�ظ��A��v��%�
L��Ȱ7��Z��rKrJ��ʙ��S����V�M�ځk*XsT$�R�w��,,�r�B���gI�-��jx���x���Fə�v�sS}ˍ ��Y�~�u����k &�L XX�3��
1���U�]����D�/7rʛ��S��,}	4�I��.���?�`�8�_v��)�e#UG�~�'T�Q^�����$��`3k(�tR��~I�l��:/�"�^T�Z���:Y�?P��0&�&�f�v���,��hJ1 �K;�Z�O�käZ1O�PF�n��I�����I��R��M x	��Ջ�T�R���睞�x�{�/�z��+�����Yu�� Ny��, (�y��$�ʦ��!&�G�E4�4��D8|�]+߱grLB�c�A�\*�~���Ym�{���gz�7b Qf298E��_V?R92U�*����ް���)�e	M;�ĸ���LU��Z�h��.x4��i�/4m����=���6����	�1�A��� s���K^~���g68��>a\�V|�k����Z��
K�����2�X=�'�������jU��&�n"�nX�\z{A���}�@�-�%��n�o�x�G���Kc���ǰ�qE���94'f)���鹷	 ��hy	��`�$#�q�8��তm���6���<����C�~�/J�,��� ���rz��]"hf{M��>�����б��_:��NZV7o�ay�w���o��pJ��b�z2Ox^>���<�u�W�'�z SG�i+z�<9v�4{9�M���V�::d��b����`��ɏQ]Ǻ/�r�C�O3�� ��Drm�
�'C��WKzNٕ\�c������;���I�d�O����k@���XI�*FD�1�`��&�/�M���W��[<�oCX��b8� 8˴|���֖���c�����櫏����L��zZvOd�Ծ<��kݦ���)��(zj�B��O[��^E�&�Қ~c�fz4�A�,w&��6c$��κ��w��=ᩄj3?�GkN��lvQޏx��<|�z>������E���}�B�&4S5�%�m����T�;�7<�X���&dY���O�@wg�HyyQ�NĒ�z"0��8يj��i��7��7�.X��p���ɚ��{�����0P��CZRA2~�E���1����H#�˭���|ۺ��W��֎h�'E4�@Ӽ"]��X��m��w�8�|am�Gإ8q�&�߈�0�1��3�#�|�R��Do }�����⿒,>���I|}s�^�Qq=q>dϐf宾W'ʕ�1WaT,�n^��oIQ����b�n6l(C�?ⅿ^�R�z����X���V��9癯]�~�����Zi�1*8|X�urއo�GaGa]�/_��N�2$���0��б������1�����x�>l�,dd�KN���{��w�*A��e/��(��_2̎y�5;&08�d���|؎�S��	Ω[-��̿u�gqQeH����Y��������R���>F�0U� ��>W,j~=Kؔx��B+�o:��0�<%ׅ�>��'�?;���X>��4s�0�#hrn��]����'�uԢ�	
S���:|������m[-���!.:�(�|��V#��L}�R���,L�%������%�B�G.��aѦD���P��J�sL�-~`��oS�T��(Go���G����5>3�؞�ڱ<�����(�f7<e����IA�V̹	 �g����y玘�ﺓK�%׏��*ދa���Y�	v��k��%-�N�_�9���e�^�\}Y�)R���g��J+�Rh� u�Ŵj�hf�̇���Z� BݒD�`�%l�wcز���pl�ڂ!zs�P��f�L�Z�"�'�(�����f�l2����$�p����z��՞�(�0?�X������H0xi �fx���Ł:g}����(��
�/���|,9�+�*Vgr���R�̑fJ�����8a�\�6��H�
 X��[������б5}�B�$�;����qGh��V��x�Q\�c([S���)뵘 ���FG�%�a= �+t�p��
�;^Q8g9Pi&�	���E����� �����Er�CL��X�?f��ď/��ަ�t�����Z!�p(R3$�ʜ0=��G�rC�CВء���\젱�s��[����۱%�M$��^Һg�m��j���'JM�˾Q�2̡�ʏe�>�$�0�U�te����^�p׮�C;J~�kY��d�A��O�a��v�ڽ�^(��4{�'��jZ�oAp�.|^�zF�<(�*{u�[Lv�40IQY���n���P�i']%RĪ�y���uLZ� ��[�F�.\���3�*�H��0a� q����µ�VG�AZg "����`b�m�F^6U:�Ҿ�L�qH^{>�{�4��+��B�vv.*sY-�T�_�e;�]1Y�f��4kje�c;'Lq���0�j�,J/(�+f`|�d����xT��75�f^�Z��=�8��ac�t���i�(�F�g�ۅ�tD���I4�5�e퓸�h(�-�`+��H)�<a�!�	��h��Ͳ{��>w���h���d�[N�0�&@�<��2��o�̵�<����y�Y�gh�����ͱH14���r�E�c㜾m&�6���Ԧ�G=��ey	nx�`wI91���,�o�a^�%}�zF�F)��_h�,k��l=���ݝ7]8����S�?jw�S��9aQ���2P�-�38l��Q��c��꩐��%G�L� ��n�
��G�%K��yw.�^B(�l'�ӏK?Y� ���N�um̮��Cag�M�-@B�E5��5|ɠ�r���tZؓ�d瑴z-H����*�GY$%�4�~����C���P��1Dr+�%;xzKe�'J&+�֠��Iji��D�9�m�>�t��#�R���f�qB)�W(Px1ץk�� �m�+	��T����:�i"��R���u�X��#��[��!��כ�bز,3�Z��CAY��yBC���m	��PRTn���������=#E!��j�$#�r���;�bUr�$!���X�f��W�<�m(P�ۀT~7a:����pL�����_8�I>�$�>���-W�����cKT>:a9�42��2E��%dPBy)�"؉��uA�Lv�H�P`EP�o��>>_�ҩ�k#�^,��D�
�_�LA�6z���R�j��f�,W�q/gͫ)K��=ͯ�.�3fLuP�Q����>O�W�������0���}q� ^k,���S �L^�٧a���qp�TN���΋���.���$���X���bu��\no>#	�Cj�����E����Bg�N\���DoJ�d3v�w�	O��8^  ���p�g��5+T:��0���޵��̻g�v�6?��Oe�c�5����X�n�b���$���O�)�{B�!s���ҏ�BQG����8b��=�X�jb$��K�;�/57����WJm��P|�ă��E�e�����vp���<���bJPT����H�{,���{)����W︿���!��',}������7u����>7�4�o!;]�@�k3��F�)�����7v�A���!
?M����Bܜ��3q}A^.��}#����g^P ۀ���oMUZ��K\�	B¯��WL�Trk�$�.�H�E��|����^��/��EqВ>�lI���	�����=s�.�;@j��b�ϝ����`oՖ��J�=����0P}���;���T��.���=��b0��8y2Ԝ4��[G�eE�ުb�5=$�xvz8H���5�i�+O��;�tP�̠��W=����Vn Nw�ǚ:�ؕi�%�zAcc���vF�j����м�L�Z�}`64�8>�q����K��D[7���������ֻ�0r���>"H���"b��)W��,]���Ͱ�?V����d&j[o����S�{B�87�񤫚��7�UVE�[x�7�a�d�PL���Ƙ�C� �i��nM����8��G�󔬳ō���a~��$��W�'�Q�Mߝ�|��l%!/>�z?k\g�+R��O��
j�Z�W�␓ڪY�)`�iZ`Q��xv����Zy+�9��Q�)�;�o�Nv�,ŧ� _�X"^�nWs��޵ݔn�����ȼV���t����]}8Q�j 0b��p~�eO�Ǿ�`w�[����C������,�[n��?��#�4ɟ9�zD�K��ц�tW�Ns�+����g�TE�O��	Pwۅ�8R����^���'!Z�z
�$�k]��zMZ�^꬙���6�[��6��\n����*�tV��A�����]�@)��~�+���z_�6m-���Kz�x���a��E�M �$Z���T
H/��Ѭ-��/�]�f�m믈
�M�l�9�6�0�d��du��$�Rl��J�)��#����S4�Z%m�۳v������r��;���9�Hl�E�@�XI
��#�3eK&C{8�q -�{�峊�
J���K@�ԓvc]�F��l��ln��'U7�x=��j��� Gi|-ob@�c1���p�]H�i��eJ\<�8U��m��E�Ɂ�p���(*f���r�Z�˭]6�@iTN��bbD��{�&ڦ�|�tia���U�����oV'�P���F0Z���s̮����e�1O���#},/��� �٪i��ˍI��;2_�+�����蘶a��.�C.�(�wUʻbb���{LL�Gv�H.���9}qְ���s��V�8�ÿ.���å�p��Yu��D0�-���̆�t�u%*#�{��o�X,d͆A
��g�'�fO�(�聴/��R8�6��n��7�����PL>���dbu=�L���ߞUj�s-' P�ZWS��Ju�l��b��p2�"XS?.��Q%3�F����W |ٱ�HAw;�۱Pdw㐽rb�*,_�p[,V�$��{�F"Q���m��=��5�L����:����QP���`8��b��i���:)� �3ӏ:ZD��`Q�+��I�mf?�Bf�@��w�s�Or5��#��kZ�����h�6��|hT]Z��� x����t̉1	"� [��yP�M"�&�_*Z�cK��5v�\�'��h��|˴��U���d���� �5{�ɥ��)�c|�c��C��vMr-
��@gA�cv�0u�'g�"�x��t7*m/�W*9�_[�sE��T�����|yIJ�Q�G}fVI������7�LL�nKs��f>\��LD�-�KM����Uv�y�6Mi�<��q�C�.*r3��S��r.����1�gryKU�Eh�H�8-�Je��[0|u�9C���"�U�*���}9*���7>fh��p�*�^���k�L/�qy�ܒ7���̻���nQ%%�Ǡ���da*��k�0�˫��7�S��TƱ#��GM���4���*�@1fx��J�"���e��0�M
d΃��'2�;j�3=1EDݾF�+��3"��y�R��ɥt�p�1��(�p�=�֦`�f-e� 7Z/�+y�X{�è���D��S6�Y���k��O#��s4d�qL�$�s�d���m�D��
��E��	<��mrϷK��R�(/����%�� HZmK@M]W�K1�e�:)c�]^�NN��
�*��Iҵb��T�沨ɥ���������x$�ѹҋ?����w��:oWt��22:R� e�$�m��,+'�"^A�p��O���U������HF�zyv6�2M{��6U)Kw7l���ħj� 
=�Ys	� �rE��)����l�y�ƀ��5&_�����hF^�KI�0��m��M=_Ȼ��Y��,(2�%�م�Q�\�J0��:�0}�vatu�tk���%�0Ȓ3�f�,�	��j&�lտ�^P4"�����%�%-��<D���Z��l�vo�O�#����qК@��^�_	�7:�=�ײ�xܦ�=ĭ� >�QH�m1�p��~��,]�N{�e9B�}"?e}�>C��Z�Ϙ��s�b`E����}Eupg�!*b�'��� �������U�Ye�����|�+83��	�:R=o�q ���X��]e(?v=�h�g}��.��K.��Ԏ�<:�U�j ��d�f&������J����Z^��<�Sh�C'n�'!$c�{�N�FI4�Q����T�^pF�g�b�w}�i�:�"Z4��.,M}6A�.�t�c%hS��`O�{f�s<���,��R7p����M���'�C�ɛ�ܻJ*�{� ��=�t]�~�]j����s�`Ծ�(��Ut(��g������
�s�*}��IJ���G%��J�{6���;��b�l���KoA��TTl '�M#)��ܗ��$5��C�z�$�hY�Ҷ���l������C��ʕ��k𾌢��åy�J�l ���Tu-x�c�$̈� T�iG��t��)>�R�c�n�l����;����a�Q����߿���鯱m�ӂ�Ʊ"!���c,����\�[�K9z/Jr���Ѧvy�?�bi��	�Le_�,b���bƐ�9��OqF^p>�M� GCY�.�R�k|�Q�������i^�A���{�Q�=����������uxk�&ƀ8��`�S!-�>���_x�j�4��� f6�|�aUi9 ]-��Q0<�C���F��$^-�⓱)�8� =��7�fI�v��tzeQy_b�EW���/M�6�pr�Ё���9�I��l!�o�]���o�����U>~8�y���p�����M��ڗ�S��ѳ��O~��/=��P��09:�Q���pk}8��ʓ:�i��h
7z��]� ��eLr���2��1��-*2��gEQ����&t��b�ɒ�)������9�lK�|d��=y�a�i�x�|Y�W�BȆ�k���*���l|;����-$f���X��n�;���վ-��j,���N�	7M;�44LqFr�>�"z�ZH�'��tˏ��>d�N[�`W�4���YT�a�_v�Y_�D�U�'��P{�ԫ8�z��W.˅�X4ĦP�etI����� �_��}k��S���ޠ��f�|b���D�;дǁ��	����.|���f�dEuo�Cbfɪ�4/��Kb������ %X�^�Q��qZ�d�n]K��Q��'*��Xxs����_�m�S����Z����[�=�搒�gQo�Srx³d�3�Bޟ�k�IL"�PZ��/�j��c����a�HJ*��x����1�&:�	��L@ ��մA�65�S, -֥v��ЖX
2�<x��[ɺ��@�m���vd�`����e�^��_˜�@��0���$f.`������sW�'�<~zN��,�{*?Ո2�|��J-]*���]8.[�'#����
)�MH�A�N�Y6�SAy�e�P�\xȵ��JkWSY'���u�=7+�ɋ>=	��Â��.}zw�SQ�h�{�fL�(�G�q���0�K�k㉫�~D�0�z&�w��0�N����Rr�];1���$�:ƼJ��E2�KqRk
�"�ą���L�bN�'��(�f�V��f! �+M-�Y']�/?V_�X]�RH�_^k�R��5��$�����,u�]0g�X���Dk�S)�;>? 3�$���l$��g��G�(ɽ����R�A�|����#o��ǐ`��M�+x$��́F7٦�j�d��O�*���wO�����a56�dG��-*�	w�'���#Xgg��AK�����?�)��"/pW&� ��_D�㨝/!�s|��o22�s;u�LZ��O�-A窷}Z�u�_ �[�����]U�~�w�&�/~�����<����U�P���Bن�o�CU�N0�J�1��Z�����w���S(u��4��v+��S�r��p�����j���epl;���5T�m�
X�x��i�"�p|=0��A����5Dg�J�Ћ`�h�`������l3�[a�$sI���3�\�r_�m_��hN
���s��l	�+3�Ts��]�$���jW4��郙�b�%�y��i���mM��z�k��З��n�faJ�+��b7�p�Gmٚ���E�I#�{��T��轧�<q�AD�)��r夈��tt����g�K��G$�Z<���`�Po�P�s�T��|�y�3���$��	Ŭ[|�������ZX,1q 6ġ\��?��/���4�m�Tj���=��ju��TM��wJǇ�0��=�C�X�3���j������Bl�
��b�H�ʵ������͒5%Q54�����5�4��9�.�{�-w�z��Zװ�C��&�����Id�4~*{�r�&}]�暨z�i4�k�E�	��L�$*od\�_��'��%����;��l��O�T&�����1t�s�
�8i��?ȏ���hL �+I��=���
׃�����g����k㡆���?ѳ�{+�����br	�'�ɯ�ر�_'+�n����4����h`G��G�U?���+���H�k��	�
�,�1�H�)6�^�����-όD���՟����g��ā*Yd+��U��7E����J����9C )�	1�%%�U{\���_�kR-�s�X��w���֣x��#�3�s@�:����!�5��T
��t8fJ$)�����f��������(f2bZ�m7�se���ʬ���]��&7�Dt~�{A�x����H;Yk{����f�'�2���%Q�[.(�Ps)� �z���\GËm�I�H��r�g/#�#�H��IG=��_&��AҌ�̂H�[<^t�I2��rc%�qk#�݄ h�;�y8�K/��:���~+m�(�uEF���L5�Q0�L�~K�'��]�V�B߁�Il��x���HV�3qG�Z�s{�S>7!&�)�X�#�W��^�]7z�z���{����^u�B�iF�n��ݜS�|�q!Ö�*�"1��t�4�(H|1�9)&�'��tN�S�:��iga�=��O��2����W� h�4���, �e@os�l�}al	�T�L���`#�
b�yI:���22��%\�����763���~��H��vȎ�c�m�~��Dp���[���8=�?kq�R=0V�ݧ7� 0*2̡��Pݹ����V���s�t����3<+"#��ҴYm��mؠ��5�\?\�z�:���ܫr�#�n�(�=��k{��������D\��)��2���7��P'��a(�	�'Ǩ�ύXo�)/ �v�ܒ�^��fj���𼰫32jЇ�c��6�,� 2-g>T�/,ץ5U���ق8��E�)d+��/�J��{:��;4�~Z���قb8�e;x�H��	��g;z�ݑ��9-��V���*�[F�K�o��!Y��v�9�9 }���򢻪�x��$F�Mc��+��n��\���[���9~Te5�W��3�\n^�fb��Ϸ9vl;�L
���<Eې�Q[?���ח$�UR�u��9�:����¿�kc5o��^uE��&p� �J��Ԛ��T�V��:��c� C�E�a,Cr_��*|A�)��������7���2b�v\TH�_��~����]r��*P��Ir<.K5%R�*=��n�م[���y��Y�Ru��'��ژ�򌡴��J`����"1�,xW�G"�|4q�D�NDAۓZ��9�;��>ϛ?�#�-1�_�a�b�;�i����-����ʏ�<����E`��[Lr�-$ma���?�$�pY�|Ȫ�w�t��k�WO]����e�ȧr�6�Yun}g�=E�s	�U�z��OQ&.�+������s��?�1�ԭ���X�$��8�k��H/��a1\���4���x���\���������w%w} Z�T�"7U�;�6����Vp����J�>{2 ��� ��q�,�
�T�O^�Th
�1aI��J�Ǎ�������&��իΎ*R�C���چ_�N�h۝�Ѝ}�/��I'�f��=��6wb�$ĕ=CXR"����X<��3�8���� ��<�d7��z`����U�Nbf<��s����t;����u�`��qB���:�D�*2�+�tK�?ٽ�`z���d}2ǀ�}Y�T�v�� -
:�����V���c:��iZ�WG��w�S����pY��`W�o����>K�d�&k6�Y���]���A$���"�&G֤7�7�� �]=�j���I�[����gzЛ��j�\f���}�!~U��
��V�'�5��и��:��1O*)T�����D ���7ǰr�����U�$8J�X5s�:;MS�.�1��z�aJ���z.����-�
�9�*wv�©��J���_�o�w�]4+��	mz�����X�AW���A��ioX�X&�B��Cڂ:q�*9�Π��*��Z�GɑˇSP �2/�xV�%!f�~`Gi$��M9b07:ۃ�����x��d���mV�U�1��g\��kϺ�vt�v~����_!�=��Ү}Ud�}�yz��)*'A&Y�%����9)�*�� $ט^l1cQg���eh}�b)��v����H&h�^y�.sfūY_My��^n���ෂ}y/ 
ߊ�2�����F�B�1�/>��nILA��)ciY�/�$;@Y�Kr]Χ�6N'�_|pq!�HY(��2f�a)bta���F�)+p��&�M��8���"��$�0����R���SCl��Њ�[Q�.��[���L��v��N!LF/�u^W��m�8` �m�Գ�f]:s�|n'$%j��v���S֍�[��)�;yWRś]�`�i�� "$�ӆ�<�Ym�:�@�= ߭>\44?���S�I~�����۠��>�K���������Go�`�UϮ���u����'��^�@*�h3屫Q`��51g�=5�Q� $"٩�����A�.��{~�30�V�V��i����s�,2Y/�h$�!�շq�o���K՗���b<Mν�!�M���v��XU2m��H�ʶHc�n�|�⠍Z�E����y�0w�8*��\6��m�0�T3e����R�����E;X�GH�b^�į�V��,6\6��8n1X\*���.K�朸Y�	T�`t���3(�@��2��^�E��׿{��e�����ew���B�4��݁�/���u�����ak��)[���\�qJfJ�,�N��X28�c۹h��R�����<����u7(5�uI����^,��"�tpcǫ���.̯��]i�Ȑ�6�&wŅ�C�����h��ܪ�ȏ�9��5�Ä
�����ɗ���W�I�<�ͼ�O#�NU�5����潕!�1$�u�j�r_k1���'��V�g-��@�D�}�2��GƵ�?^f*B�kW���B^�U��!�"�+�����ZLi:U�"��тN:~�eaQ����pW�ۄ���қ�[H�K߅��r�S^Z~��,[��N��:�Ӵ���ة&ڍ�k�q9���ԫ�L�
�e��P�+52=��;�D�y�S]�?>P>C��^�wߗ�w,����b��t>q!t=y^FνSӔ\�hC�� �!�U�J)�׹���"S̘�Dx�?.�_c�0�� |R�q��h�����ZV_^8	c!hB� Q���h��3b c%���s(HT����{��n��De�N_����|���}����d�]krg�9��
�]�)]�س���U��@�����{#�O���ٸx����S3����c����Z��ss�����s��=MԌ8
�H=�彫��.���_�aǖ����Й�JT���T�]���<p�u�������%�= ��l<�hL7��QEl��!����H����֙���aΠnB*�������'�aX���-R�.5�]�ܭ�����Р�
�8=�*��ڝ�R��E8"�M���Q���@ӽ���Q}8��ڱ����>Z�G>��`ʍV�H��5�N��+��5�<�V���[�o��~6x��-P��'����iW�>P�)Q��3Vmq�����x�\���]�W%�j�N���R�|�sR���|����K�1���B����EbN�����>��ۡEo�i�1���L&���˶ٟ�ùcB9�]��b��mn�K(޻U���*��`��+��[)!�K����wP�v}��7��k����|�R#�*-S!�7m����~�0�i0C���73��"�B~�d8�%IT	�l\M �Ҫ�	����2w*��`�J��SE�1�z���)�ME����\0��4�Na?�-�㏝�5����L����H ��cdi>�B/��p�{�fΘ|��dɪjI���[}(���.���y���,ﷰ	��SD1�Mv�#������5�U��T�e��j2+��k�%]K�����ilW)7$�'��.\���:��+"��|I��@�[�ן�`�:��Y)��ƾ�,3�%�!~#�*�|+�~��.�>�I�[����Y��ǎ����`��&�[�Z��d*.&�X���r=��M.��%��Nɷ$� ���$7)�������=���+�0 �c�аIZ-��mRn�mcG� �Z!�b�
2},Ґ���L(�|��@P<��ar��{��t�nt�c����}�������_g�F���p�?WaԆ:��Y��g�f�V�,6ٓ}( Ѳ�)�|:�@��"�%a_�Z�ƫ�ק'ÏP��/K�[<[c,��t>�u�ǉҡ6�Fw��R,*�%��5+�悵�i�Ƥ�����3L�xhE�3v�]�m?CqT�P���h�Q���Hl\�P����'�LGI�����d�P j8w�օ���b~���`�t����`���$����Lc\{�Q��x�4�-�
+D�>Tq�(K��c��w�B����јt�.$-.�d��D��a@ל�\�P�pOb|��`��u�X��-Vf��,q6 Wɹ�f2�@����1j��A}|GרI`ȷ,��Xq`W��"6{߿����Ha'6O�Q#%�	�7#r�5�AK��n:��i2B����3���"(jTZ~ԋ|(ӗnr�8��D�y��_�����eI�=t��Bo�Wt�2H�k���)�Mk�{�J� �iwѸZ�s�9Y%}I��v=�MA�j3	�s�p�( �<Ll[�iU�<��f�B��a0j�����%C��k�^�}�o�i�y-��(x��+C���p��u�r�ɗY�ܚ�oc��f�%��P{�4X�.Yl�S�����"��%�?a�h�Y�ZO�ϧv���X�x$Lh����K���Q��\���3*�e��k�6�M�#�-���  op�"G�vZt�pW��sA�}-�F��xt���'���<Y�W�SF�v�=�P̍���f�O��$��Fi���x��`uU���=���Z�$qk�2Ķy)�ŉRV>ַ��X�����F�5������0G��V'DxEB��,?��[BT4D���]_��{d��=�*�0� ~EJ�%�+�j���D��R��s� �֎�Lv�(�ɤ�� @G�繁���~����a9�%
������ϭb\�MZ@�3y�4�d���2�
݅M�-y�j���)��f+�r�n1E�b�:��C#P��-'�qͣ�ag�3�#Ǒ�z3K�3��(���g"�ݔsׇ^$Y���2���;uf١rJǯ4D���֘�:N�3�����ȰˑY��(y�}ȅ��*E~m�˯��u��{	|lFMz~��Pj������{T+[Mh���m��f�5�-���:gr]|�l�o�l�7H�y�²әN�B݊��5~D��.���Ԙ�Y�%����w��K��o74�2�Yh�1P1��aF�!��!7���l�)�}|Y_	\Zp�KK�����QB��,����'��L�0m�ʵ�}����pb擵�L�'��s�$�dulbIg�_@Qc�)�ٌ;�(��q:38�U%>ͭ���Vƍg�ᾒ�Vzca���NK��]���>��m.f��h�Fq��d��g} k������\]�m@%)�������ai�8�ΈK�r7���'M<{W�i�*�k�������L����rHfü��3��ӥ�3ebW�Fdq�X��Xa�G��tM��Pм��0�!P��Ψ_��h�
~�x����H���˽t��c��ڻa�z
H���"E�y�����k�/ʯ���pA�����;�q��^^�Sz�@����B\ާEvܔT��P��fj���������KS'Q�|�w#.���s�n�_�����I�� L�t٤���xWb�7�y��x�8�5]�� 	�U>@���U����tϓ���:�m=b0VX���h	*��٣+s�rD#�&��s�6���U�L�l褤��N�3�S6q��l�Z1�$��C�ʯ+�Pf�t�'g,�|q��\0�������?��ZB�d�����Z?��\�x�G`GC~���B坦">i�`�aR�V%�(H�'��/ �e%����$��ó�8�Yy(na�*t���Z�H(�R	ѻ<�u�����3��Ȯ�f�w���_/~�I_�Px
f���9>L�9q�O�"�)5h�f���2��dΞ+bN�B�6`^�	�N/ި�A�����67T�*�` ^n��Y�T��I�)�R�9�ެn�2�BJ�)jk��J�u�[��dG�"r�gn��㼡���RQ3��KN��l�^@�P�-:	��oӅǬ�	M���������ӏ 9�u�\��0���|E(%5��??��M'�� ���}�����nt"N$A�h���>XܭY��ߤ��Y[%�VM�� �o~v����X���.���dZGW��7Ē<��f`y�d�����p��\S�N��\�oP4j�3�VEF��9_�gJ�.�{'�[%Q0����t����yҹ�jR!�j���[x��K��*Gb 4�U������z�~��)P,���K+q!@x�=/\�h��D'_�700����}�m 3�������R�=�$�3Kd�EU��#P\�t��n}/��?�y����j��Ͱe��e���T�#a��:�G9�Z8���K��Y��]l�J0V���xp�����Dh�K��^Ү���L�_�呍WO#�1���c�4���N�wɣ�BT��^��~Q�a�N	;ۼ^�����=]hl>!g�m��,K����,�'��CK�P�Ԧ]�v���7{j�P��z����6�G�� �.��݆x�G.�+��V���{��P�a��&j���{KܽF�=JK�Lш��a��v��$��WT4�r`�E9��H���K�ʲ��ϑ|���wI�󙖅p<hJ���  iѳU�AJ;��Q'�$a�C��;��(w;�9������k���q�^6�}���~.>�����Z����c�`ݘ%�s�:0��W
�2SZkEZ��_5
1�Z؝� �
b�����"�:�$��X-���ܧ�����x���H���^�ƫ��o�#� s)��������OL��B�oXE�0}2�e��덴����R�F��z���/.�O�~P�3JA�/�wb��-0<��a�K�b��ݳ� ���@=O���T�P�����'=�5����)q�bh���X_�]A9G�Z"s�߲lkL��O9	>M)�D: Ho�X��*��G����uE�H ��|=Q������'�SBJ�����|�9���S�ɨϾu�/�~ܦo����5����0���(3z�l�=��+%u-]��n��kR���A��8�t95f��.>�u�Q!���Go/Y�ؼ�'��_c&m�ˢ�t
2�;4�+gj�iĂF�K���ha���C7YL���~������~L�e��MK/�c���ir����k�� m)���9u6m�i��$C����/���H��$J<~���vG��0�G�'���䒀��!����m{�#z<���;§��3N^~���-����\6ɏJ�~�m������L�;�*�\Yw�5ܿi�G냹u�QI��X�ko���I�l�>
��\��z�y�68*�T�c�l�.+�đ��o%0o
�e`�-N������=�z��Rg�2h��Vd���ΠXh��z;�&_���oqI&�U#��\u/�N��a�Fh�)��~7u��2Z�Ԫ�&d��&lcy��?�3q����[8ne\���=�۩Ӽ�h��.�ܽdW���Wc^!6��1��A5�^w�����U�aL�ɳPx���o��c%礗j�o��4j�܈B�9�VK祛^������$�P��a/�b7=Q1�sU���L�~&:�ħS�5�����$���ep���K�d��6Xm��H5�����OzO���@s����;�s���J��­
T���F���g�	,�!h<C���
��r��O�+ц�Pz4eYX���IJ7[�o���5,m���X��pے��`E��c��V��8���@%o�~�o�dB�m�P�9e�uӹEY�Hɂ6�^4	���4�5�������^g��ID���KK�"�-;��F����-�V0�S���nT���v����S���c���0[�l��N��ȧ�~?)��J�K�,�: DO������v�����֟��YJ�����z�=�#b������#���=�0��j0t����GҍD����"l�W��O�X��d�+��G�?[�г�z����Dp��D�yʑ�%���oPl]P��v��k���+yTh}h����7�Clh�Ak�>l��̅*;g��9���Q@#5����B�R� ��qCa�ՠ�j�ھ'�f�Сs��b-�n�(��S�f�ȟp٠= ;T�)aCŁ'E�'r?v0>�;Ё(C"]�r���,�L�Q�h����h�jG�z��Y�GD��߯X@u��ғ�R_l�a�N��Rs!��A�ͳ���|��X.��%��9*d#Q��i*"��JT�h?Ǉ�!&�/5��
,���1o�	�`$O�݊�����ޠ��:ѯ�̃Kb��>�D�?9�h�@�Q"��9m� K"Z>�<��1��O�Q�SC�Y�;O�#���b@bN�]H��H�uIN�����PF-t.' �,�jv YV��#����G��_�A��)NolNP�nϩ|#2���3!)U��&r���<e#f���Y�;�zFk�Qpw���T(��]n�2F��D����X�Hf�=��g�YE<��B��}��'�rXغ�`Oj�<�^�h���*�T|���y�D����N ����������i�G�hȭ<��5$ C��&U�c�s �*8�p���<�ϼKD�8S�).c�˵ٔ��D0` ���p�K�0�Z�p�1�	���,>Yt�k���_ηz_�w�FM��'{�����:ɣ��(v��ɪQ�����w�L��w���$Q:���	��HH���0&�����=T��7)^��TNDk�>G��4N���@6����Y��h*y�q�hp����ڕɏn�^E�m���bF��>Q��]��[Y��v	�,>/PmR*���]3�[��1��¢Y�ͤ�����l�`�!�H�0c��S�.$�k�
1�ӯ�������n�����Iʦ�nM嬺�!HJt�hs�g?�N;����l�D�<h[$�%Sσ��B��0���r��2���ڷ�Ϭr2~��[�"bW���
�_e�0��%���%�c���x��ږ�u�{kƯ��`S�3��H3���;
l�j�(��.��1<i�V�]1�ݛ T|��^X�x�V�y�$����$����r���4B�N�C�J�"��(0M�GH�f�(;�OW�Q��T�R����Q��-B���u�֢e=�	�N��]R��Zʙ�
tU��:�XЬ�CeNԸ̟N�|P�OC�Wao�}v_����_��Y������R��n�>9��0���������3T=������]ݷiV���20,��$��?�<0J�P?�*��0!�������ӈ<��'�V.?:���-*�C���u�<�%�A�õ��I�x�Z#9X�NF�렣6�&�Ղ~����a��E-��~����R_C�_�u�l�,nJ>bZ�q-�w�Q��O���ؚK���T:3n��*�9���$���:l'�v[;��>�] �V����L} 4�`�v�f��x��/�W7��X���+=Y]��wI�� _{���x>j�r�h1����l�K����/��EL7�o�e��^kO�E���1��_��<���>P� �����B�2t�������� �� �]�1�@685_��3��:U�[�\0�cZ¬Zb�e��<Õ^*��ZZa�~Pab�cw��`)�䄏�9u��X��V�ro& ���S�<'O|" ��~i���#��U~���E\佔{U���>&Fm���'������[� �z)�|C' ����]N�(6���B��l�����ֽ�p+ i~��f�c�_ST�p��~���1f���=FTeY'� Dgs�n\��YUB#��L9�m�1��uv��|��7��62�<��,T[r�SE-�O���<m��Ϛ��2%�͎2A�z�4��L!�߹�u��M��z�=��:V�^�X��[��ST��^Bm����?�� �tk�q�p���A�<?g�x�����3t?�V�Ym� ;E��m����X4Ģ��5�\T�G�N_"Pĵ���N�`���0mv)�҂�
��k0l���)K����-�3־Ğ��zH"5X�i�p�c��-IEe�8~k5W�t����H��z aȡ��sOF�2�K�]�Z7<���֔5��m����Xzn/���à����F4UHO�8s��<(^I��&"�?�yu�bq��sw�	���$9�և�`Q�ąa�Q#a��M���\�꾷jBs�O���S��y�4V�������X��b�V��������9�����~�obr����Cؚv`���2۳���d�=&�,��m��ٔN4AW�q��H��-)��o��{;����]d���P���24���k�eoEk�$:/I׊5E^ ��W���s���wu%T�KS�\n�^�Rc�'�$�� t��C��Z��򝦛V�1z�4ܥ�e
���ת�Q��o���8/mO��|�����_��5�1��kX��_���
�.PS�h�Z��p)�b��O�lpN������q�r�Aqp��|���T�.�n���T��ɀ_p��o��O)������e|���~�ROZ���J��!
a;����%ſx��������P��6�J�g�#��+vJ�(*�5#a%���{z�PBѷ��������jƏ�u��ז��pD��/Iq����ku�]^�����?a��Qan�<"
��K1����dgS�_[{��ٿP�}��HX+��i�*jH�jD���b�]h�w������������=�L�=2�4�*��)�W8̽�6�?G�:�V���rbD�R,ZP{~M�U[W=Pau)��zN5gQ`�L��>�p�QTϘ]�Hf<�W�&h�*�L���J�����Vg�}���I�,�!<45�/.02�u��^�� Z��?�Y1!�T�.(�c�B2A�*Ɂ��E+��ы1?Y�~yu #v[� �Ax�zw�b`|�b��n���e��1Lj������S9����s,e|VB�WCL`.�H�15���>h��'��u!��el��o��7�l$"��X�u,E)ӯ�dK�a���V(�#��,f���`^��5�v��>�U׀,�P��\��tu�_M����"�=]�X��}𤒾�vO�p�<�WR��V,���r���a�=}��.R}�$���u�f&���Y��.*�����#�Gw�<��S�Q�S�y쭉?�-p'�驔����E��������9����������޾Hf���\��kc���������Y�L?�����ZZ�N��|=bZgU���5+�u;ce
��8��%	=5�9cԅ���IUS�Sb;��
�yWN`���G��^m����	�n�]'Y�(�$�%	��~&�IӸ@���j-����L�� �|;���%_}~�;��X��qb�F��b�_wi�skw�7�a���ё&�+�2�z9��ŧmo�#h�����Rz#���i"��?��@�J����H+$9����a��X͠�O/shv@�]�u�3��F�\��M��j7�e�<y��̧��=4)�ԚXIQaJp��t�xdd%��GW�O�1/��B8�_7��&��H[����[@fY�� ��T�۷3�������@�V}s���vI7��yv;��37}�6Ā��ŬO�I�>XԂYX���Q6�K�x%DƯey(������ '�K���3*�o��90��'��z>��:b���<WZ\G�.��g�ܿs��'E��̋�rK.�2
s�-���p�-�}�6V0q�E���qj�н�KE���BX����p���L+�n'-�s�{ ��b�%��{w��������o�(�n���z|���`�Z�~��!P_|o�3��:��@Ո5���)��_#*�ͧg�'$;��-�Za�� K���{u�����ܓ�r�v}���}�t�hr��'E(O�@ۘ9m8��r+�Dh$�5R�No/k/L�6Zi��o�E�#	+�㉪wE�X��짟��ԮG�x ^����>FM��� ����/�O���9C�|]�`��y'���r7��+5k����!�*�d��+��7��@n���C4�ˢ��k1�ː�/���5������7.��s~�"e��8i�B������,@F��ɑO7�{����w}�#{F�9���|*�@�C��A�����2H��ƽ�x��%ބt�697N�S�R>�z��~�3�@������1ҝ�/�L�,^��Y��J:r�$2R PCQ���"�e�=�9"@��/�-�px���V����;���3|�2���-i�%ľ���A?2��n7�ߵx^(`�z�X*��̎�Q�%;;%���)�[����#�s�.�]�%�� �ϛtlZ���;����aIeK(l�@]�)�՜�\��Q��!�Ih*�6g��nq�ے�?�:�3�
�A&����"ᘰ��Zx�#K����,ēZ�;9y�, oK2��"?�w�<��}�96�Wdl����[&Q��5~�MyH��L�a'�gq(�.�2��/�)��f.��\R����:�zW�-v��+w�+��Cg#\�{g��s�<1)O�#Ϩ@TV5[�����FY{%��:��Z��t��O{�_�sq�w`)��tb��#_��b��1��	1���q��������#E��w3�0������]�Ia��M�u
�rhv�^�&�i���jBi;�BܻH�8�v�\�Ӄv�<:�����\&�<���=N\�)ki䪄��Z5�� ߼�������^����֥���/Õ��&�Fn��qQP6�m����@�1.�1G��3V̹���}� ^����u�߰����.MV���[/�,���83�nY�!����\U;�/�8�y@pb3uC�A�:�������f���Q� ʷ|*�*�Э)=8L���ұ[��:����/�����(w]�y�
� �;�y��'�u��?<�=2�i}Tf	@���a����\Y6��Z����>>[lW�fx�/¸ (*�u;ڧ���[&�#��m�p}g�����I��U�Qm�o��k�r�OO%hd#�)]�ϥ]�e��6.�|��RK�?��y��>�R�SMMؼ�9Fw�^l)/�8���HsM ���\X�n>e��h��us���6��V�Y~�].�	��KL��Z�0Ha�p,mW���}K*�c��Dh8m��y��|6V���TfT~l�y]U*�zq�x��2�aԸ���k�J���9EE�w��V�w?�V��|rخ�-;�gc{*l�\?ڀ"N貘���=/�q'� ���if"m�|��@��|��ސ�Zv�H�G���.�b�ͅ�
C}��?>w��>�=Tv V>-�Ӥ��-÷ģE��/~Sx�"x1w)֕���!�jNv5߁(�w>��(\�9�"�t$��� �	Wg�����č�$��$��_Z��/-��az�B5������h���ű1lt���8���>}JgHb�OF×����%q�$�Ch�1jv�U��GNe"�V���6m���>K0��3�>�o1���MN��C���:���sQXȂ��W��}颤���Mq��L沼�B��њ*�f#��
����V ��#���z������ ��e&�\\:Y&qɖ��i&  m�jXg��Q�K���ЙL�KC3����3���JS��_�T7!�����>��wHn�mO��t�>"�����C��R	�ӹ���M��~�SC�y�ـ������r-�7XY��,cWtG�tT�U�/N3k�8��r�X�Ri�L�#9�@6���#�K�YV3k�De�߁ă����X �_f��ؓ���|�r�J}��e�k,k ���,6�h��^լ�;v30���ۿ:�g1dq��Ƞ�&G�7�Y�|=Vێ��m�E~�_.i�T���j&��Y6Syd��F��5��I֪o&�6:�,w�(������ݡ{�H,��'��)ͣƛy�fzR�{Ï����a=i�;E.�<�G?{.�?Ys�(����uB��@��]�OR��;��Υ4}��-y4ٺ� ���һVn\{:PԴ�d��+~�A�S���N~x�Hlʳq��5[�j��=��o��u�����75`��@�m̥�����O �������W��|Qo1ņH�BE�Z1�Sf�(��tY��/A̬�3q�74{$�۝M�*`�$��cx�$�eW��Ni椛�Ӗ��>�������q]9��v�V�m�з�ݚז9=ns;��|Ok�I������)4�n���s�UQo� �j�j�i�7U&��dݣF{��a��#��p���L��0���c���Z�:�����
��}��f�o5��n�I�!4G�r����뛧Q���,���i�5j.bL����E���4��Х��>�Kۨ��8C��឵M��	��6��D?J�1 ��*�j������U㸎P2�<ܬv����s�/�������}z���No�%�FQ�N��A�=�ڶD����p�kG����]�O�����fX{��g�7h�aS�v�Nnw��'ԬQ�nv*�|ֳ���Yl���F��0���֮5�L��sg��R�~�<�����s����g�c�s{]��X��h�Ģ
����GkS���1MhY���M�Ҥ�1��.��@�K�EW�0�D�e����"�1�����8h6$FDu����	AFP���j��8��(<
)�J����/���i�sK�飍\������6������V
�LV���u5k?�0D/uo�*��q[-�[K a��q�ώq�;�\�\w�R�B���J7��g;�
�(��2\[r�/�,�pi���BS�z�2��%"N7����Vh����Ƹv���0p��>�ѓ8��Q|i}�G�������fW��g4�.G᫪+�����4�o��G.�CE˧1P3!M���P��*,�?��MvT�o�Izu��lf8�MMr���V�~���f�V�<�������K�ٛ$���B����g�y@�i6�蓒R�)R�P<��?�����9��z(ͫ���{�Aެ��qVFb<�bv
HA��-������ٸ�b�����6^�V�K�`��/���b�<��:%�8�"�SFc�X��w@QT.,�(�cX���,��ڹ[|�g� ���E^�s̅p.;��SGf.f+�qR���?deL-���Q\[Y/&�� ��žD�f���e�f��TwXO�~Ѽ	j$��~x�8$M�;��~�뤹	��vM��ѻ���Mw������X�Q�p���vC &�]��#F���d܊q.�R��C�MȻ��m��f��*��ZQd���4�IZD2,B,�A��������g#��t��-�HWS�sR< R<�w�%�ߴMZ蚙��b����y�_�,ѡ�>i�EW��8A�Q(~���˅J� u� +�e٘[pT���V�G�lkm�R�p y����i�����iv2��u2i�򔁸�$���:qZwj%G��!*m��+����/�ϝv]�h�����pE@�vGK�G��V�.����7�.�H�Pߠdq��/�ODܓfV'W���n=˫�43�b$��:�C�y5A8�@��!�컥-o��Ϩ�.z
��:2���8�B���SX�������D$~*♘s�p;C<��]"�B`Na�2*j`)N����<��/���l�Dh,/�)�o��K��z!a�j�>�Y�r��$�W������|��=��Kp��:�i��0����3�EaK�EJ~$w� � }+5u�+x�:���K����.�I�G";���_�iV��M<6�q�����`&�T `lPj�����%����a�3�9��	�J�;���!׆ш�{ͣ�>L�+4��^}Aop���`&x#���!@wm��.��o��!˼ >��
m�$<�lQp�mG2&#�����,�/�� �S��!(^h�J�
d�]�uL,w��Ά�m.�`��^�=q_�h1v�Ao���#;rsm���<f�1(Y�J�����/vfGS��&�&� �М�>��\�� ��ݱ\=ZZ ��E؈�}=^U�u������o~	��<E� ̓0�� ����������!j�Hɭ?�:jK�z
���ۜ8Kh(�qpΐ|<V��Ȝ]2��>b�_!�����d���[�yk�,�.�#�F��L��ޑ<�a�s�[K���zEQ��Jb��ܶ����v��IEn57}g%Kc�5��ML��h��`�݉j61YJ}Y�R��^�MW�eq��]'�g�:�\(�"}����B�CE��C�S���b��7��Ɇ~/�3�&�f��OzZm�ٺRl���$z(�3=��u�pkd��|�5X@�Vm#.��rY!�����\}pn�M�씒u�E;�����W�g�D�{`2Η�\�Fq��R���I��o4:;�ޤі��_ϑ��x�4v�߄�_n�j3z����P"�vj/�#���Ϯ͔~������%R�RsC�^qu��#5͙�y��\a���fŵ4v��h�J���Q ���zz��iM��ɛ�=h��T<B��LB��"6'�ѧc(�R���)z��"��K�&�qF�-d����DF��L���.�tr��A�(;(@�l矠h � �g1+o�kE����%&�qkb�ƶ"=	��wQٍ�c�MG&)NO�S�=̝�w&��m^G����H\R\ 2ڂp{�>a�$�nP��9�#,Y���J��K�Z6�S�UJ�v[Ӕ����q_im�	�+B�ѫ�n�+��n�Нqu� ���0
!u�"|A�3F>t��ӌw��,���x�T3���>�qL�rл�r(�Ύ���g�~�rf���-���\�x�u�*��#f:�>��X��d̉=?i�I�6M�ż��`��ȉ�D��nV�i1��yǢ��SNd>��t,n]|\�'d�e���B� q��&��rѢ �⯙a;��2�=v��FE�%e=y�։�Ǉ��F'V��׹ġv^:i0؏3�eg��r�?e�����u���V�'7Mg'W���/j;�h�"F���EP�Q6�0(��s��.�����SL���b��#tb>�1�o}�\�N����|Ŗ�A�DRB����C�H��p��#>ok�h�g{-��.,O"1�ѤکV�o.�o"=���B�pO.k�N�<B�#����Y�o�����enP������5h�L;
�C,����y(7,d-�d�)��jD�s�L����T��0iр,R��Xҡ��;�qpB5:�~ZJ}�KCG1����A"5�*�K����Pm��H��<�΁������k�и��w�j�А�Qx�Zz`�"��m���n3s>_�Qs���(�Xeojx�CfH	M!޹N��XʫV^^�^2@F}�-H��������_��o@%Q��x]��W}����W%��H y�gu܅��Nk�e[�Z��@]�CXx�~��M-�,�"��_l
t�EL@�l���R� M~�N�����X�[A�!�v)�-����K��fT�^��dHi �v&%l��*l���ϖ1��hB��oB�5P+zţ�7��CJ�s�{:����¦�\u�!gզ���/�#ny�{�aM��D���⽸Hyq��saޔ\�3�x�G�!*��\��k
�(�U��k+����j�a$s|~��^�R[��˜���
�݉�ȕ��ߨ�7��s؈�V�<����>^�RoT�8OJ��_��X��')�V&=gܽ:�.�έNɜ�B�_�pm)B��)D,�2�=zß���q�M�H�>����}��Ϡm�JB����Y�+�9���o*�({#ϣ\
�.��8�����\����_�+ð�j�"�Mv���A����җ�N�$T�%g����d��ʁ��P��T]g9]A�0��������N�,d���PA�W�J����u*�;Q�������ˈк��1f��t�^�~"cc#ph!�x�H4)�	�9tfbԮ�[J9��l�5��p_*�Dm}�[=Z<��f�N� �.9�R�T�* n�/'ORl�ά���G�1����:�ZcB��'5�����y�(-��&s}��_J0)���g^�A�.88�b7V^�ÎC#V�CԤ�$�-7�l�޻�}��f�6���	��&ǖ��'�<���8}ڰ�v{!�<c�����P��?u���\�X�5���ȔX[��Ⳝ��|��B7��o|���F�1N?y��߂-�.�s#D������%+�4V�0\���Z)�C\k�cqvm\�����[!�/]���jd��wc!G��� r��>K(������?+/XD�y6;�&�B��Y����͉~l,&��Vhs�������,fǧ�dX��C6��TJg<J��	{�Ob��	G4�{nؤv�nT��Q��<�aT� ��Vͼ��l;�n�Ct���J�Zb�^�T�;$B��4U@�i�����~2�F�Cs�_�݋��O�F�PSǌ��r�>�� &q���Q1ڬή��+C��X�q��kьa�����r2�X�-�x�[����rS�P�I=?
χ~ϗn�s�kҊ(�Ӡ=� !��#��5��JBϸ�Kp�u�К��H���R��?��	�U��w\��M�iBW��r8v�����v�ی
�r�g0�@z3e t�y�[�5�k���)Mݞ�������5�y�,x0���1�>��e_�%!I�] 2)9Mr�nեu-W�&�XI�iԴ�M����;��Ʋc�h�C����a�;�v+��]0aW+Gn�^uf���������4�MC��e4��`=׆@����k�\���Ƒ�`�b�V�_���O�>ŕՀw��b�U�,Ư=��b��-a��G��Sjl�#r��X����%	Q�Ϸ!��v�d���^&���4O���%�P���C�k?��BM��hD�X����ǌԃ�#XG�Q��|�"v�}���O�L R8�j���FX�/%��D7uMW����"]�E|�݉��3K�,"/�s�:�o�Gᅚ�ӚXr�F�&�bs2��y�ߕ�ȗ�1����:+�u� �D�F�US������e�J�!(���Q�U�G;$y�W�U��dA?3P��m��Q��q���*���b(g�N=�}���&(���yS��K]��Km���Xs��j��F���Z?�{�sU������o=�޺Es�+o��>�Mp{�w �r�9��'sEtL��*�TV�x�rP�8��G��(E��y�D~���E���P�lH����+d[
ŗ�v���H�m�:L�:��lc��w�a�Q��}j�$X��{	��#\i��m�g��N_�2#�W�O憿��Ǫ�v���s&;$J罖q�_�gDzb7z�(�ʃX��_�]�d�h�6��D��F^>&��`��X��c�OM�$�@aP�����1� ʘ-����-�]^=³vY����Y����;�@C3L� 2�@��!���Bl94�����9���,��Y��}������Iǳ�mԳ�L�2�����Ln&���3�*�G--X�S6]�~t��d�g@t�X���t|��쵪PZ�6�%# ?�0�g������+D�R���9{O):r�f~��������Z�G]k���&W�����l2]��������ޞħ���H���h�>J|`@��^�"jR�쁅��C\�В<9ƹ>Q�����U��\�DE�->�㥦��d�e��Lm��+�VS�� V�_�:��R>�Ώ�O �ο�jO��b��7m�<-�,��R������U����m|��e�/�Յ�Ϫ�_�(������(zwPK�Za�W���(���=�&{�;�r��:�N��YI�5�[������'Xa����*��I����w�8V�N�<��q��$E��aW�Pc��Ie���� ��h!�xb��ח�}�
����V�E̤�u
s�nj�n�oKQ�Iwb �Å���n^�����%<��/x\��w�
�O�N8�_�n�?V�"|~�Fa��;����.��*�`��x��wUW��Iз�5�$ͼ�A)X�IL5�ڠ|Tco�� G-�j��T.q�&� wjhpz3��u¿[l^��B2���,��ݤ�}�*�.�oq�t���*nr������g2x߫����193�����!6_��O��S>��R�Zq�&��)���^4DD�nMV�qD��O�˷���~`X���{�k9�G�_���	�]�%���,�(��7��'�z��Q�~�t�k��Y)��ht�ý�6��W9�ne��,�K1�p�,GH�X���q�c;�5P��43�A���IZh�,���(͛P�����і��w��x��OB������?R����D�o�_V`Fr�2y���`��;�7�7t�FV*�FG'��`��*��NQ�g��
S��\3e��D��~1�X����_�y���C����7"j�g>��_��2DܫƉiI�t�I����X�ݔI{U��h��C�zq���O�q��+!�>���v���nV�"�j��!Q4�wK Z\˖GK���j���C$��@4X��	���I>��LĸP�^j5��A�p�1�Ujס�z���únv��
֑K�Jm�߻"�3`:S���V��v%D�@[�[��J�&�#1~��,��V�n&��u�=�=Ҵ��i7�y~(,���X��$BO���~���5Řq�`Z<�� "�t�X�*�,`p8��'/e��]�����+������|H�z<��mYO<�{;��C%L��հ�R�>� n�s�$
�G [|xV��Jd|ǬX�����Ym���t��j���$�n{[$*ܗGx<��ł-�r��<��^e�����l/�8s�!~���$��N���2N���tpK+�<�0r��U�q@������r�9�?k��8�գu��U��V������E����$�r�+z؂	�B+�Iܻ�_�e(�}z)�S���q��J�����hX�5�%LNO�P�^�*v���B c5����3�Zz��q�w��É�;Ve��]S�`�.#�s)��'�v�`ʕ�Rx���G#��j�V=������ik�¬����w��Ua'������]�}�����d7����E� 7�)�C"��0dF���L�o:,�69Y ���0�心+�\�xv�y6�	�{RR����nm�-5y�3�"ӂ�)�UI2����Q�c֑��b �=�*t"�ޮ`U�^5��Y�o/�ʇ���$�������S���F�m
�4�rk�g�o�mr�h����W<������At����L� !����h�W.�F��hc�q�,�%��]��:��xP�7�&��S�d��̍����=$�Ʃ�p"���jѤn�6>����)��l#��j&���T����A���4���j��$Q3�Ŝ��8��*^]�آ�
m�ɣ��K�@iI�J�0���S�S���MT�x"�{\�]5�Ν�<�ֶ\(s�1	
�ԡy.B�-�_��6JF��c��MS���l����d��9�л9��ErP"��[���lG���k/�	T�9�!si��.�����HI/'HQHC���r�-��E�35D��O���I3�� �D��o�����+Jm�e�S?������*�0I,���9���`��ObC� Mu;)1E&��/�%�~
��s6��%u)tI��rkAG>%^��?��\	[�S��{�����"ǺDx5[��3c-4���-Utag�wP���f?�PlCc�y!.�Q�,PW�(��h��p�[��t���fcc0��Q-M�f��%\Mǎh�.+��e�������h��ƨ����saY��w?�S�ն\�Ud0�\�BʎX�Λn2vt6��F�7ヵ~���ۯ��TE�7ި�a����3f,K8���Wħ��*�?+i�P���&�%����U��Dv���}n��Ö����rw0+T��DB�?���i?��թ����T甍������66Jb�Ms��4�#��k�~�&L�ju��13���,�rF$Ōq�����Z�C��Ula{��h��ːX��Z�ߖ'0|�߼�E��p���ʱ�|97?y��ŷ��Y\%� ����]s˅�LBI�S� _�O���S��W&�=b����I� wk��|��g�:YjR�
h�������H��R�E���BM� ���-?�H�5�Xy�6b�,����T؄k)����1W�lLK�z��e�S�oR���><�]������ɡA�y!$Gv���p���	a��ס��lD�$�h�k>XZ>m^-�!�����6���N3�G��ݵ�B�Iʭ�������0;�jJ@=N�����OP�;���������\É�CsG- �1�6��d��u�Kѹ�^����|�)���HI9Ȇ�X�+�s����っ]��f�l�0�!�%��h'1��jC<G�g��q'T�(O c��Xw�rbL暁#�h�ѕ�'�KOs<�AR@��?��}�������l㒲��b��Bo~6-�6	"���a�1�!�8�i3]��eH�kl>¬�Ĉ!��b(�l.�]��v�6D{����4,_�{�~9�УA&2���
H�����d'��g�'>�N��������S���ܕ�9cY9)�+��҈-�����X(�����˨���0�n�e��4 /qy�(�h����� ��N~Vf%�\hcp��:"�SC��[>,��Q�����dId�����=g6�'��#�s��2�,��]���F����$Q�(�v����<L�kef�Qױ��o�wbD�]�,+}�ɢ�,��{�oڗ�X�uBWw��1�ٴ����_�4M�2L]_�Q��=���߉㭆v��+�Nj�uP�y���wwY����lEփ\H)L�&!lso����U��?��&��,Vj��P��pq(=�7�s̺��b)�m��qpCN�ykCԽW\��im+�s��
s���pZ�7%ySjr�:(��6Djۡ1��8C.�cAT�\�E�Q�8\J���c��"��E�q���qRL:Ó�O�f�5\�왦}KQ�`}�ϫ./2�~����2�fN��F�!�Y��U�JC�k�Κհn*H���KG��<	NL</4��v�H:$W*]�'p��i��ĩV����~s�ſ=V�%j!���$ �i����t2��җ�NyX�	�z�m�{��^�=�z)�<3��͎��/`�a�-	���pr24)���� ܡ&�9�y��H4gW׼��u4JvA i�P�,0��C���A�����~>9��om�%�~N�+���y�_lT�x:��&2�q����v���b�lQ�$�8
-#/��"�"z3�	��+�t�cQ��~J"��$�!"F�=k%��j�B����T�U������P�פT'��q��ׁ������m)B���%i9G�l)g�Z�_Ac"zJ���Z�hS�����Rz�:~��/9ddN�.�OT�O�~��N���s/����E�������ܘG��c�~aƎoָQ�,II�;v�)�k6�;\�z�gp�_�o�X��Y�-��BI������"�+�r�"������$jVV��Ol���̗�a��=i����[?�μ��1��;XuoTE�����)����U��d<ֶ��w�� ��,�����0�E�����M*\x�eK̴usV����Jƕ�h�{iU[��"Y��2�+ �@V��H9Oʏ��]�.h|�ҥ���֭�w/�&��>s��+��~r˥��KMʨ���y��cd;�`˔�[>�#��e�/���i���'I��g��jH�һ��| ��"<����>J9��9\����ڝ��w(ل��g�4,������^&��]�a�ɽ�1�8 ��l��H2s
�ܧ�3/�hK.b����[���̼�Y>X�Ƿ���@��Z_��?�����؞����֠y�o�m��S�Qً�\���"΄�[�X{�hk�D0!��|z�Ew1�8^j&��j�O��O�����s`W���1���~nZ�@�~�d�Β�GN-JkH= �A�+�MP��!��6�����8GZ���-A*	oe`�8���z׹�Z��ˀ�ڗ�Xb[B�I7���%�l@��v���I�?�%�T�H}��9X7�q�y��0qg�S~��>h�1����\�Nz.�Z��\J��t$[����,��̍g�c�1z�rf�1te6���J)݁�%�X\llZ�;�Aj�ӽu��3�c��"J��+w��~n�ᜍ��ч1E�)�f�0�j��^�!��1�C��KTk�6�?�d�b���kՕoR����~��)
?<�W������Y���$�4��Q�l�u�|e#�YYY�w�u�����20~�6+���x)�i�����p�!���KZ�0$�~�p�M�A��8�������.�1?bW�9r���ig���G�HL�p���BE��Q9��5V~�3�l>� )J���q��3z�$�����,~ˠ��H�wFӃ�� �ⷑ,4�^B�7�������2���)�CU���Uq�p���0N���T[�g��S�o_�?늅�5�Kv���Jլ�%���p��do�!�cJ�f�Gh��#��OCȣ�e����h��f�m��t��~ѩB6Jzy���c
�I< ���(S�_�����fu��h��yK��.���@b�5�'��`��g4NB>�F�-#AxxU�F��g�M�2n	� �wӕ��7�Ek����w��W:�N-��uqĿC��~�\j~���&�w)$yF+����2������@~	,t;�F��h�����Y��*��6�iu�+��?g#�������}40Lz�o��$؁��}�~Dļc����y'�*���n&/`�ZM�<�\�)\2�O�N/�&U���,;Rˣ���r��bU��*�f���+�j>��4�0�n�*[���Ԁ�������0���CX�d%�s�M]��!&}�7����6�V��t~���+�EO��򿹯+R��8� ���5�Q�>��|ߋ���O�\��Dr�_Zk0Tj��YȦ�PU ���7����'&u��tL�����.��c�h���	��4#���BR��#qhЍ�p��h&	�0�$��?�l@����fk/��0Cu��F�|֬�حcʨ̽-����[=k�h�
�� �V@ ����r�gUӴ잳 ����Mb���*xr��
�DӪ�\�.�jٟ�T6!*-�&��=���a~t�G/�	h��ة&:%Q�T,	�t�^���fSBi�E��U��Qs�~M6�9L7����)���Q���{J(BE�a��ӗJ�ū�
��$d �\���4?�,���
�L"��>ԩ�z�@�B7��GU���}.%s�=��3?ZS�̙jN�ɠ\�/\l�H�?�Ӈt��N�����xi��z�=�g"gb���/���V�h�x�74_e8�9�.�V��-q����'�l���Io���=� ����������Q�<o5��r�ΡTMΚlkЋ$�Z�#�#&����g��J�ա��Rj��P�%E��B�ůǷs٠'�m!�6Y|�7Mn�p����'�A�M�պJ��ݝ���ڷKn�i%�V�ᦲ�-�k�@�fDF�r;��V'��%I����7���+��:��%�f�x��kBp���Yi��=������=d�q�����Ĩ�^�Φ�,`���V�Ȗ��Gx�kV{���y�[�t��7A��[�J,�R�t�m�&Y.�q/a�1��M�-�"�A=����w��ۯ����������%#?��~�	15z��;�qRZ����&�Ɯզ���vq�w��jn��1�����2�ǝ��D���T�xv��Ւ�GC"Ft��A�("��χ���n���1���$6�;?([���1��EE$(��F��OR��h"��:�����R������yl�����N�s�����S#:��*Qby}��<uT�6.9�8�X��QiI�����f*^�
�R����hZ¢��$V痰f��+������ݲqj ix\m���\%�^9T^hgsEO��7�6�����8~�WX
ڕT�����,f������١4�I���n�Ijq#n�a����^L��n/�$���j,��-A|t�W�9��,X�9�m�N��/r2�[P���m�l��beNǌK� OR$Z��5x�c����Җ�z~�JA�C���X1c���0�(w�*v�e��ĝ5���̦��=H��X���_�@��ڍ�(�$�mK�p% �}�J�= "�#,_܎����y�K�Z�X�V����h�FzՎ�s�o9�����o��ޒD4�\�/G�P~�}eU��8J�1R�n"���"����7�<?��k�=�����;�����>��x���(���{G908X�\�����&S�ř�#q����i�}���ZQ���_Tōt��� w��#RO?�jӉV�}
�;��n��J�O��/6沟gD��]%]��w� �w�ѿ~��m9��]J.���Vd�?�����3�_�]�q��?a>�n �%3.��^��e ��?@��3��H/�Ҵ��yE�%�]��/B�8�. <Cҧ�ғ-���#ע���`�)���ד�{b���H�.P�9�3 k��H��;,����r�H���h�d�c����/i��
����ډ�{E#�}C(�+�5="�t��1�e���g%Gւ�WG�zJ�jS�� �a��&E3��t�bR���[dB���3	��m�T_��>ɄӾw��GF'_o�����"�Y\�-ӑ��K��p�}E������f�e2[ Œ�����A�T�!l�.ڔ_�aU,���la)+�.!����L� �C9V�Vm�էW�D X#�>y �g+-N�^�E)}-U��5wO-�����Z�Ѱ�DE���$���_���yil�Рz!%R�=M����5�(C߆8���m��e��n�UI�y5vrQ���^)�*���S`�4C2��ߤ�p_묝BqE~P �j�\�]�I����s����HES�ʝђ�͚$�j\��B0By@���l��ۨ	h2M�A��k���o_mZ*�$���/O>�v�>E�f�Fo�M�����Eپ�`^};�I�2A��F��"�')��/d�y�_���r�\@�x"a)����8<�/���&W}�dL�ed�˶v'�P��n����h��M��(Bf��%/��`j0�b�����B�Rq�3L�0���6��<5O��˺p�(C/*���{ ����L0��I�qW��Aw���n4+��۫�U-���8e��E��8?����Pk��10妝��ȕ��bէ�Q8��7�N�1���l��枨�L�v�iU�VT����C`ch�.�p3�ݚJ0�+,c򦴔�vaX؅�?+	꧅���D��l?=Ӟ��4!e��]S�� �+E�%Ca�gB�|�P�?�X��^H�aa;���p���b'�=��z�F^L#&�����p U19�	.��Hb���X��du��־��[�1tl0���LP�����CA������lV�'r<��X���lE^�����a��0��Q��//�����D�wG8\��ii��7e�(J�Um�o����ɶ�����s\s�/$T _װ�n	�Z��:x{"�,B�� -o;HND�>n�8��M3���SC�����S��,+�4�v�����U�����)B���'N,{[x�K�o�W���ZK�O�2��Glʧ��<y�-�=�5SɴO�$��(�!*bď4v���g��j��k���[iƾ��8U��,�N��t�
X�(1]��r`���bR?�k�"�(U��,| TK�76ק��X��]�%��a�����)����2��z�d�b��YA�g*Et���bI��}���`��{$7�[�W�Fwl���)����TQ�TP$�܅b8�+5�E
Y�"
�Z��:�қ9cI���ԛ`z�1��Ā7�������̾>�T��޲Ab�Y��>'�]af�9]Yr`�V����� ��d$/~U[o�yV�N�ԝXN��gs��	�Z �u��,�9=��U�����Ҟr�e�`	\�9Bbd��f��|d�"���m#v�Fw���_u���^�z�R��(_應��LP{e���<�|�����`��	1�Ů��(	��%��6��9}v%�q(�3��n���]I�k#���rS0��L�W�'Pxs�������E��P������NZ}Da+!�8���$)��йo��;Ao��*g���H�7�%d���c��E����6�1��Vئnw�t�'�4F�f�b�K�>�w���X��^fN�T���!�
�kp�7w%�E�O�;��$�<I�e�w��E�<i�	��-E��J���h�B�sy] Ծ���EeN�C��JŢ�eSdP����!_��%W;���0;�ǂnCӊ��{�e�D���#���ig:��@:HOcKp1l^�~@e�ϕ���.����^���Ӥy3���H�P����!�Σ�^��+�.K�%�g��wB�[�׵g8k����!��Ǿ��Qp��A�'3T��E�Z�q�D�8c���u8*X~z҇irK�(=����
R[�r���7�����,D�l�@MC{N1��.�)2�����e�\�	Iќ�A�ON�8�f�M{_�*̊�w�L�n)8�2[�N�r1e�[�3���ƪo486x"��dz�O�(d�6�V�i�[�FqE�Ox^l�1����:C6u{9��w>BL�w;yχ���'���Y��Ɏ��©ms�ج<_����"M��dm�@=������p�g?��^���OV�_�,y�r�	"�y�}�����^��m#)m�^N����5�YRx�߃�zQ�/�L>x7�_��̕4~���Tx���iX*��ErJ����8�C�WL<Fj�&"�k�D �2�Яh{�s�/��+ �P{�x�%yq���Q�װ�&�*�mi6@"m��kO?n�N΄FM0s���S(ۼ�c��rv`ms���_ԕ��,8��a��T��̝��ԫ�����#��Zi᪵g��D�O�]���lف/?@h'0-)�QA|4�A,�I�`�ę���֍F�g9��,m-��R�-@���-�K�T���]3PJKT;$�q��qh����JD�r!�W��i��Vef���Ϋ�xIuqD��99T�=�ʹ��:�ŉ��-V'G�\N,:~���9`�ȍ�[�������2Qq9l�<
v��ݩu�2�o������W��y����{��'P��i��&�Pԅ���TW�ܓ�l_����_BQ�S��}J'�Gp�������Йj�7�d!V{��Vrv�>�Ct�����D�����
���<�V��Gv�5�����Ysr���z�
5|�<:�>���0Hr;z�Bhv��A�tp`��'��kEn�`�T�r7#Z�Oƚ�|'ɜx���$=��4�� f�, ��b�]@B��b�K@������R`��>5��0��A���"$����#�ʝ	�9�%�,K�d�$������7�U�Iq���?�}L(;�.�'��5����r&�B﫢����f��|v�p�~p������x�+�Üzݖ��UN�e$
ٸN`sL����ʍ�A`�L�#���q0�� �k��=@�$���+ � �zftd�(��M�Q�sx:dU���,�+��s�p]5΀
-�m�|�@"f4*!�YĂ�H�k|@H.�f���^��@%:��^k�� ��D�p��`�� g�[���M���?E����?�>��M�+L �b9p�ѯ8����2�+�7=Y�*RPW���2�L�����.~��o���c^-~�%�{�ENDV�U+����i-Q�1Eq�ޡ��S����	6��T_�����n�s�i�I14#\�鵹�ޙ�w�'�� Ƅ%B.Ksԙ��ؼ������I/]�XC�����;Yy��*aE�^Q����-t��Cw���=�b;;�OE/����p�I�
\2����\��zK7���}�k![�h��1h���G�����s��+C1e���j��K���2�<�o74K\`�}
6-�Y��)�FuK��Xr+rumT�W�;�O}H���������Q���<�͟;��+K�9�p�֥���������~���]�B����;@ж
�,�Q��*E����9�XaO�T^�}tAM��0��Y��(�g;�M��ȴ�s�FZ��d�<X�)r��m���B���e��Ϭı� d��-OwY�Z��_�F���5�����h�V9O��Τ�a��w�"�.�����T�_�-��0���q�5�Zc�}SG~�M��l\O�����?�N�h�i_��:����i7�0p�y��V�_��L�f������S�Z1�
��b�L�<���Z?����~�pRQ-�E���b�w�����;E���&r �oE{
�C��X�e�j��1��:�tg���V���R8�X�{ve*�z�sC���F�c�k��x�[}�@ˆ���Ҿ�d#Z2�����5�Qw�-4|���W߈��I� L��M=��+��+����XZ�B��a�U
؟����~����yB��щ�@����s�b1P�0�+0�V'�A�A��lsW�cn�j*>B�8!9�E�R��H��Pt������p�������#F"Q�ْ1ɶ����}�8�q�y�֩���(�f-�^4�����ޡ3����mm1�IP4n7�*�is?<��-%�i?�yC��*0,[�?~L\5XQ��$x�ǵ~3P壑(��y��:,���D�
[L'�Q��b,�j�k�9ʹ
{����n���d��N'�����znJ5�\��<{_���	A��K�K̸+�5�8�'جoFxl����P�rǬ�=^���Po�Z���r⨒sJ#�q޵��L�C|p�]�|c���	*��������To$LG�Mi�Ĳp���4B�ҹe�K#I���������!�F�A�?��$�m�:-x2��m����u#�Bz�q"�S�37�S;����x��%���G�E�-�͚��s?ₙ�RVr��-7;�k��(��j.�q]�������^Ҝ�2P�e?0�ѨJ4C�F'�V�i̵΁�^�n��H�vb�D�G�R��f�xN�U�Q� "N�S����xʵHHAal���� �d�}�i�>"� � S	�F7$Ob�7�2�}s�e�}���옉��%?�2e�4�+u�Ą'
]�#��+*IO���'��NbZ`��`*���6�=��K���jʴ�h3#� �9Q�4\zI'��Q{1��	��1w�$hA#!D��Bҫxh��;�,���v���-Ԁʖ
�ӷ�bU���|�}h�ua�%�䳥�;�L�"����+�S�Pys�o۵�f�*j�#W�^�}���C�+���3/!�5�΢�(���Rނ����h�I��D˵�?�^��] m�C3�����7H7�
I/a�K��1����|���N�(�����9gt�Ђ�i	��'x�[��koK����ȉ�uP��}�����R���-���t~�X8RH,훖�u�6]���{J�A5j�����>VQH�>V(=�z^B��s��F����N��L��Y�QL�������t]��4Z�0��Iѵ1!��F�ADr�=͕�j%�&�U>�.p��;W�目�U#	��H�|� �H9a^bt�kHjf�d@��0��Y�
��#LT��n�.�yr�cG�Ky�:AM��cN�D Bi��܀F`��{�J�?��&M6˯
v��{����h%G���i�U���b3����	��c+���y����i0N<����vΐ�K)�TK6NYnp���>|>v��X�K,�/NY�d\G�Z�B�V_��,KT�!_s������y�� 嵀��7�?k�5{�t�fO��d���D,�	S]ձ���R���o�T3l�Gǝ%U������mݣ�E�#䥿�P�Y�&�8�Vh@#��&s��0}�o.�H��R)��tuN�׼y�X&mjs��5 ��:�2u�����+��W�`Q���@Y����4�� ]u���B:���LH�%�%P��9��luAS�O͙��,�����!��$ń^@��Z��:f�i�J�,o����Z�fy|i2��s��T@�Ͻ�	����Y���!���J����v��I����E�VNJ���M�,�5o�@e%��!M��i#	�~S���z�d��,���|�3�m��յ��kT����,���s.��>��@�(m�)���A�0P�-A�JXe�ĐÜV�l5!;���G�a	o
����_Y��[J�S�C���_��)�n�3�Ӟ�f���ۏ���R��:��q�;�W�j�٦��kyo�E;{�����-Q��H��ܼC�f���j�3�����W3y���iD������7��_�Bj�O���.O]�N�<e��	���=����fdC�yye��,{R��gM�FW���vK[��-�?dh3���S6A+��F���0ݛc�I�p��=W��ɱ�]{�7��W��z��%�N�����z9w>�Ͻ�p&����2r��ZU��"�x�@��D�0��n��#.���� �q�*��*�G�(2��9E@� �&��J�`!��/ɒ��h
iY;ܘY!�3�}��~.s��,sN��|#�>��L&3��JZ��2j�{�p�1<����XwPl1�g"o�f��օ��\=Zm�
& ?�Yp�n�]�ޤ%W��n�ҷ�*�F_r� ❪Bk[}M�K��(TD;�Dw���xMY)}�xLJ���tX��%'�5A��~�O[`mzaɰ���g��bvsp�ӳDMb����dn�X�m~����7�g[��p����:�X�_��I�s���(�؛�/<�dx�EM7r���	@1p�<�F,(�#y�y��9-.����_���J�3��y$����Zq����h��0�h1�~�c��@�޸5{��҃������c,Y� [��vwHZ�%��G������S�d_U���?T$�N^��pF [cb�NY:^*݃ԏ���֛��8��N����d`�oLL����S/��^����6:��G�S`:�8!�K���O��S,-�[�<y��ZM�>
�P�|���v~��Qů�L�N�p�t����ϞG�ιt����b�uR��~oJ�t�p�-U*�a�����cW���sz��TC6�[��H�{/?�.�c�� ���8�?�D6򋿢�ľ��صB�/�����sc3�
���H�>*��2m�_�Cf�$�D�}���0>3袪�3>jT��s@K��$�Dy<�����X���kF1j�Q'����D�F/q˩�aq��~@eJ�����	�&���G�)�ͷ�h�V��,S��/���9_]��c�Gk�ᰫ�I`�I^n�,�qh����~0rh1�'���X�G�W���si<�LX~���xL����7���q2��k�d�)�d����Oe���*X��A�Um��ܿ�?��t�p��ռ�<��>j�%e�3�p(jhj����4ms�}�$T6����rx�*�Z��C�s�����cj��9���VCy�f&�*�X�0HɆ0�c�
p�����.y8�ޝz�}��$��hv�>ƐBy3�	� ��� ?ܬ�T�;BĔ��V4���W(���c�d�]����r�y�kx*V��W�����~5�o��,\��g����g�a�e����垈�m���q��0!doR�sb���L�
�c/�0	4"Cب^�p���\iV��D��Oec?�����P��n'��{C����ǃ�:r���a bw���
�b�X�.�~��[u��j�Ab�'t��� ����5�LE�jt�53q�eӁXaU\ΑW�e�"�����(����k��D[-\Cl#����C]"�wթox˪����S��F�5U畽�:�$L��.+ЩL��i��k�y�R��K�6��:�d�������(O_�B�ٳ6A�`���f��g�m��B<����N��/`Y�^E�>�XGO;8=l�tD����C䑍 is�o�|�k�d��P�G� A�d�峀4'4O�@���0�����1�5���ݢ~���t��� ���(+��
�0�a�C�/S��QH�x��^	���.>�"�Q��\h�]�c��|�\vtv;_�D̪���D6gI�-�m4�"�R�?`_"S��gAڱ������pW�8EA�j0�3wN6�/�f��9��B��Z�W�Mn[�F����53}n�)����'��4�Gh�� �3����9*�7?{]�%.5����dT�6z���v'{�:��4�N�~\����;�r�ӢS���V*ލӥ��3�J�־'s��ysD:�M"�����j�{hR4-�sÌ�N������؁��t�

oG��/� D�~6T=t�gp-����olT�8J�M��I󔼓����>t_[�EXK#��Nb�jvxD����Z�g�2�e�*��^��k'�T��Vօ�Ǆ�#�'��˕M�� �%���1�8�i��8�N�fS����^�	���l�K]���֏�G��Bڳ�d�_o����X�5I�4i@Vn��sxJ�]�ݐ�S�����<�4��e�Y94��`��(�>'��a�0��
:�p��'s��4��"*��`c��K/�8��K^^r��@�P�~	���f��x��C]���.<�#��2ɾy�� �><��H����Jm.�h󉣲<O�Фc��G��?5��҇i��߾���(.I�~X������v:�I�@��Z�g�� �rx"|�`9�}m�@||�p�cK��
ܭ@�p=��#4j0�L�◩#�(�wiDuN�QѼ"���*��kօ����R�S'c��޿gC* ��'e��B"�ݢ	�ѫ

�x�Z�j����PZ�y�bZV��	�%�:|<R�J��'��/:��T|�ɤ�v,��Q���#R-<�s>�<�*�\gxM#3D�p�;4�'T3�QA>! ������G�:b�U��ɰ�GtZ.:�.��s�\'�b�����.�4�����
�3����9��v6�˸��[t�6��U�@���6#����PxH�ˮ���)>��h�X�����IД� �x̮̕����D���L�&;� ��&3�&����҆~�1�8���y4f��9Dֶߡ��E����_�BϿ��x�bS�<枏��:'�0$�A�C��Ө��;��8�ߴ=��R̐4��3���bD��ڸ���r�l�C��O�X�E�?���x9�3v^Y��L�y�Ĳ9����|�6qn<Z���C�-�H����>�]���O`�ځr�OxY`8x��9�̿�����(.�9f.2���>E���1�I�_�L1�����ė�T �ҕ�<�
�k��n���v�-��:�u83C:Z��w�5��[H�#��zʔ6�P,(hr�@ �̿�y��a[@�J�z?�9���o~,��B��g�F�.���aW)������Cm�^�n��O����v�M�5,0_����KH�b}Ve���B�8<�&{l�fؾL!��E��7f�@-�ǋD慐$[$|fC�5��.� ���e�mpʱ/�<���s���SRfǊU_x����y�^�	�@�Z�!oc��W��Wx����
�o�Ձ��N%P�?K�6@�8K�o^P}���|#@vT�M�������_i��hS�ɝ�{�7��g�۲gz�B�$sJ�˴Z���[��u�����(w�j�2/�*{�S�����1m+��.������K�]����Bwu�w��y-������l$�r����%q�T��=�|�҅-o#O/�p�&L��c0<����^�\����>�Jur��u6��Ϩ�ֳ%� e�v�QL{�����!	�ϓ_�Zo���*�<�mɎ����U?͖;�H�?���@����tpWG�	���-U&���Bs�������S�v�\�1R�kTzsӅ.�Si��!<��Ŕ`�`à�兴%GO������sQ)p�����7�֓t3J��:q�q�KR�ӬH=K�Z�7s�Juݠ�t	���.��#�ɣ��ZU����v�]m�m��[�/�e��oR��1t)P�����XoyC_[�2�(*�Rn!�P!�#LK��?��Ǿ6L/��K!kP�:0n�s�U_CL6��g9�HJ���I��2S��y��] �0~O𛗶�9�Z��
I��{��V�,�l�#�?�~�K-d���.��Q�c�����;�p�����ه/r�R� a#ݦ&��$�a>�p4�缍�$/��^a�!eT�iLJ��i?�\Y�9MFP^{��4�5JT��sW��}1�����vw��m$hg�l�E/	d�m��T{7+�d�gE��`K��͂�%���H��6��2��ĉq�$_��� ����pӲ,),�mܗ������oQI���
�é��#��X�1E�sk���i�xw=!��\�0��ؑY�pLj5j�e�i�w��@�Jh�(��1BÏ�Q���2؇�x��b���T.�xk:����q
xe�o��g�{Ҽ�R!l�y�N�V�s��%p��JE|�֙.(9d: �!� �ѐ/I?�۷���2�b8,�c�â ���E�_BYJ�)�����.�
�ɗ�)�ڤ!�7���3{�ɴ��^��t9~�َ�fh���� �ް��Y���}j��I��t64Y/��7���T��7�B'�"��d�6�bRo�i{&M�`�e�k����n���n@���Mt�4�_���j�B���xǁr�$�d�<���|��t+��g�/S�63b֗��il�X{y�	r����Bb �cS��ې)�|ng��?���<��.(�-,u�<v���N�e'E�wͼ]#�$��O��
uc�iZ��}���p(���ƶ�L|�"˴3�K6,k�=��3�3}Ƀ�#?v����+0&=ƥퟯ�'�|H�i�9�����&���^>��n�ም��W� b*ep"?9�z>9N�i/���Pu�:�����Ą�����7�Ǧa���N�D���Z����Xꀺ+� �l'838'�T�	��"����Z���~fL#i�=��r��BS��5M��0���3�y�����ˤ�!&\{��$�ZaC�;R6L5�m5� ���]34oXFdlIl3�}/�n�НcQ�Kʑk�0[�>8�(
Zt}�4��������~t�}Gj��2б���a��u��3��y���J��6������TMg�g~�I�`b� <���gI+��������,�a�x��!���4n,tO�Pn��G�<�O��o��q�>��)��$��St�����I����5��W���L�3;����\��,%��K�G~�}�v��/S�i�)"�Z��WF�_n�o�;��sw�\u�b��'7Z��'��c�#��Uȓ�Sy���0I��xQ6:������Hbv�����#"���08CRE犭�0>:���f���hq[��� �;j
�a��?�ꤻ��x1w�%T,�s�f�'�ڋ���J��ߺ��U��e��8��ⷒiնQq���yPk�)~��ڱ9�v-�?��ma��4�37�&R�W'��[�Y��8W#34-��&�Aޮ�`�����tّ�h����5h�O[+�l���ׅ�rh>�M��06wI�cw�Gdӽ����	�Le�#���P�͟L���2
 �$i�M���+�M�l1���IR�{/�D^��H/�ж��mI4$鑸A�΋ڛ����eD|�3e�lgG�&����x�,�T��.�(�� ��{���!��3i�(�Z/�*U �T��[�B�'��$H�M�N�T_Xp�0�PtR@�5�H��%8?��z[�x �X��#��@���Ԯ���cG�t�N8]X�Tحr���vw�x�L2I���h��h%�������,�ĩR�-xd���Y��qWHD��+f��i������fz�L�!2U�R ��;�.��݁��Vf	����3e���x��ne�8��X��,�@���:�G�+�\���t��"@�*�w�P�G��/2=ֈq|8�e&�ȉYEڋxS	�3w����5D�تo��qw��=��?���G1���� /F!0��#�B�_wެ{�t D^iԀ���N���]b�Z���~��%9�ݖd��r��M�rYߺL�$W-\xS�Ừ�N��U��o�ڴ�2��#*�ʧ[3;��n�������VO9fH̝J[I�����-��9�;�ʇYA�$���l��~��̱A�|�-&�#a�E�)��wpĨn6�}r��F2Е
�U������	��D5����M2�����c�*������*��6=x�����O)lCj��Vޗ��\��f�B�.N�*c�K�ڏy�����+-�3>�ߠ�@���;�����p�.�j�u�h�qW:��Tn0 
N��^����T/�xy�D��Vj�2Q��}�`JR �6p�5X��0`�w�2��k�b#�l�c���m����m��_�RJnz�7s��`A�	�x��ςkK'��$Y�6��{�2�#69�kk.>�%*�!�\^B�� �ZNxS��� �4��-&�cnG�^¿��5�������K-PJ�`x$HVk��#Fx�l�q�JYz<(��A��J#��E
�k�	�d��&A��kl���6n�%��Ҫ��������"���]SiR������4o������V��ڝ��Z)'ց,f$o�i,��1	@c��P4 z�h�Xά|:*��9�"۴\c�L����@cc��t��Y���&�ѐq��ޝ�zsNf�"0ۃ�8@�:*a�
p�ce��^��`�\w��O�2x��#�K �~{�?�R��O!��h�v4�K���A�Jñt������sN��%��F/��H�PW�T���钢��D.��U��
���Ÿ9A�*-��5R#�Y� �W4k�6 �(� z���	��5�%3،;y���AU+�8��٘��cr�����(��kI_�k s�@J�]��3*�wr���
��8_v�����{i��N�k��֩%F�� �֦ŉOI?C�J8v�\ODR%���;��d����(>�Z��;WZ؞%v�s�\���pr������W�K+vͬ���ϰ� ���hMaU���=����X�eE�T����1kK���OD6�F4Jp�=�t�|�;�)������1܃c!�; `��3�Ij�+���'�
�L(6�o��厄h�H�&��;G3�[��I�$����el���~�ҒτfCK�Sh@MV�����|M�'� �|�~�����i;�mW5w�U	c���nr��׉aIԉT�>��cq�X�����7*bȦ��˕��}TK��4�er���F�M�?�g�]7~]*
�H���p8.!g��l�%�؎���ct���ڢ��+r��O�������S�������8%��-�Wɜ@:�rJ�����4&�G[�vQ�a�l~ǚ�>Ť�u�i3�U�/��Fl��U��V:��8�Im�J���%SΝ�i3hSq��0�=�Uac��̻w�;B��}�)A7�lq$�x'Rk�Z�f'1�m��@5�K	9�a(^}.�Tck�P���.(Qz��r�말	^ewY��j�`������,��I�AGJ� ��xK���I2ӥǵXrx���\�TN\������v�@<��<��&~/��e[;��hn]�)3�p�VWr@��eO@~�;a�a5�Sz%�u���J�r�N����B�SX��+-uz�(/��eeQU�~��'���G "i�$��L$R�!����%�e��������&t����ì<�2ٓ~��m��fD�����yC�W8�	�;���H37�zG=dY6e@Y������A�ѩ�Z�+C=��\���a��ߕ3v�DH���x�L��y膇��ʹ�0)�B�_B_�"��J�	YT(͹�W���7a�eCn��N�M�'�mJ3sUq��n}��"q�@�ǊJ�OP�/����'���PC�Z���Fl��H�G�Z��Т#��i�i�"".e��9pد����3��ģzM�խ�+7�����YM�8�0�|Л���
�Z!��!	y.�*n�X��m���>��Rwg�L�L�ԏHSZ,�X$��H����Z>�Y(:�J~X�\a��d�;��0{YQJ�Q)�0�O�\X�����ͧ�^<�'hE��#��鑞�r2\�*_-�6�%d�B���N��!������!���Ct��V��[	�&&]��.Ҋ��F�	K���di���i�_�(5���Ʀ���/�����Hܿ-e���'��IU	�"���[�ʫ���>�0f\�9t����P��ʱx$y�����U��$ǝޑK��@�a�[��i��0��3����}(He�,Y�A^�)�zI`�@�;��p�D'��՚8/�8�U�}���~ÿ�0/B�~G�?�]1��v����g�0<�aa$(R�U�1HZ�=k<M�o�rZ�8ͼAK:���$�FV��^bQoG�5��b���Ɋ�c�	ͨB�f�Xf�Hd��Q�"�qpDkZ�j@�ֵb�g<��� E��Mq.0�d�m��u�MЉ x�}	�F���SHIt� I�����V��H(ef�770�#���E�Ԃ�U2����)i����`f�����z�����`ߩڵ�E�6�P���/�\ �+-��S���%�=�w{�c�_����z��������b��S�T�`��f�h�9��E����cv�1g�xs��:D�ʳ���۷����+OZ;�Z%�פ�I�2UFQ���E���� l�o����zs�9��O��;)/S��F^��O�2�c��K�E,3d��b�w��*���S
�q;Ƽ%�A;'����Vr�	P� 
%nH�{�*�h"����L�2����汫/�Bj��EKW ����@l}�!��sR^��
L�[�L��9�vbk8��w�죛�5U�ڨ��@��Ȋ�%M��z��X�;K�Y�䫕��Zڴ5|<c�i`g�5�H+:���{h��'8ko^�5S����I����w��6݋H%�	�)TFW&�v�d^�/������6�U��I�Ҳ2�����i�	l��U7�z�_�w|l0�z���0!�!m�s�'�X�U�+_/���r��\cY{X�C'�P�'I�+���-9͋�g�֣
��HM=ݨp��a�\څKd����I�v��6�V�zH�$�7�ɜǌw��]�(N���2E}�[<oE���!�|�;8%~�I�JJk��n7�oވ��x7�֨wb����j�"�h�Hb�g韰��@�F	�U��%@uػ9IKNZ6�|@���9����~�zn'��Zk�d+�Q�=b׋p՜�N��552-�]hj�_�N%���ӈ�|�|J�%@��W@�.7->3���d�i���%Vn�ݶ��.�j������k���5�N�ԭvH�8������M���.i�A�:�Rj_�X衆�f��Qh���>*��:�_�&3���&!N�v1S�{J5?���!��R1�Q�	9*�U5��z�M_K~z��)w�o���ar�I_�X���-�
��!L�۫�S<_����.�J�j� �5@�[p�"���z��E�O�PQ��\>�G��Q6ӊ�d1�e��8��x�T-v��puմ9�|�-HK��/�чI�]!�����)�E������|UC��ͣ{�N��PPG�z��,Z&��e������Xe��)���~�n��
���K��4uA��H<���>k��X�n>S�7�^�����+����gQ�V�x��%>>�rۃh0��L���~y�\���mj��ԉ��=��\겜}��]@Z��7=hOQQU�$-M�V��ȁ�ij�y���}�e���xx`�����ݍ�
~���c�b`!��60s���R�(�Q�Ǌ�P)-n;h��-�u�{f�4п��=��}�o�覇-��Q���_@��O`te��7�c��K�5K`�-a!���pdFܤ��In�V�r�g��:W���b�?��l��K{���:i���"�S��/�����*&����t���h�g��FSv>u2�H}�ͭ�³�Yݳ'J(X5ߣ7Dva�����Gx��f[u:th�L�������hBX?�{�:�����<�o�n�T4tF��	���b�ۚ�r5��-�y�1Ch'Fwa��^n��_;��A�^ΠX@4��"�A+ͯe�B m��.��B��D�r�5W�Q�+�9Y=�������|Cq�9�x�S��ː+�*�Ѥ.��8l��(�mʭ�����.�-���?Q�ӛ�)�*�K/�������5�d�������4D�t@�d�c���~�g�+��{1
ظ,���41����@�P����!B�K�H�����S�3��j� O%��
­�07SSIG��$b����)����јT.v�iz�.�y�D9�zʝ����	��Z��}�G�N����A�OVj��v�h�گ!��(�ot��O?�o��6 m�Z%W ƒ/�2��dC��{0Z8���W�c�[�� 8��QJ���47L���E��
>�D	L�8K'_�N"=�j�y�Zʻ��$#�QZq1�k2�y:c�\<��5Wo�|��l�c��J^����u� Z�W�,��y��֭ؕwA���ܠ�5��b��llf�g�[�|��#�џ�*`5?=�IÈ5�6�N���N%%�ue����Q�Z�:�|e�LU�0�I��y�V�h�j媽3�i��Wߤ!RX��|^�6���Sn)��w����,�אM,Px��eSf��Ɏyv� ��e�
�M*�g��L��l���#/�s�����8�*�z4�3p��v�=i�_U0����4��m\�C��Mğ�6Shi�:떮d��2�i���x��(���|� t�
���t¤}[ ���N���i��)���H�_C�m�|��FIS"�R��.�O����U������#�u �K(�����i�֦A��X;w�39AW�E�zE	k��v��Im�^)U�\s�(<U[��a�a���[�I�p�`�ݮ-7��`�_�G����1Hʴ�H�-s5M�/�b��:�l�����`�Pi��Mr:3m���'G�F�ѕN�c;n(m��N�j7��SSo5�k�L��$;�D�V��}��r�ħ���X�p�E��;>��w�<͢I����`昹�E��$f<e���		C.\��kD��}<�cfVZ5�w���x=^�a�/G9�W��@?[E��K臥D���5i^����Fci������+
_���a�1�W!n��]���Ԧ�!�K�Z�m��tX<���o�%��_�|��sۢ?oe�b�5d�2 N�6�K;쿡�R���D��=Sv�I�Cl�7b)���_�����|5�]�K���2y[~�Ev��1�K�y�����q*�O8�]#�9��w,��^J+��[ԢL������^ܵ�E�s��b|f��#d�[��w&���0t k��7��[I
�<&��G��� ��\�mձcg��L�O�^��%؍w^b!g$�����tb�L]==W�a,3$Q�M��5�u��a�
/QVb(���'�+ڠ�֚����5�����������/I೔(�J��ѯh8�%X�1-B�Kwe��<NP| �v3���G��ճ\����ݬ�
�x�DV#u�;�w�:ռD��c	�s�#.�M{�m���n��,�+Y���r��ǝ������ѯ��xq���:��r��@�mw�� )>��ȧs�)�����Q�DI4i��Tj��-���1���H�&��
�J#ۈMH���]�I@g8Q�����y�1�)H�SFN�H��x�8G��c_��?��[��ꀢz��_OV	(��� ">���ȕ!/���>z��j{6%2Yg�rP� ���/:F�ܰRG?}�M��Ʃ0�x2|Q�'+���{�=��#��5��.�:J����s���e����yw;'8�폈�����#�7������P$u���,	�C��L�p�������5�v:��F3����^�������f�����m�j��,��@��<�E��nrg	�����w'���=�fI�LM�Ӣ����<"ċ.�i4*�;5�&����UKZ('s����K&�;�+�ԝi��N8^���Pc���w(��'𝶬F>m��������)X� T�7�ܬ�@��v��0�܎	Ǧ2XP8`�p�i=�^o�NB�YYz�ZT�ㅺ���|��K���Kȝ�6#(⅗��̕|b��Z��]-b����O)y$��DF�X�-�K���+�*@X N�n�$f��7ص/"�i��!�S7�M��xq�i{����7�e8�X��D�_����2�;�� �n��/�wߜsZd�Khժ�b���8���M#��g�<B�͢b*��&���L�ưVX�-�(��M:��36^̩,���+����C�}�'��W|OD]@Ӫ ��A���ߧr���N��MЧ�����Dg���<�ȺMb��x���@�#��*���Qo�n�D�ՖX�r�n�,q�:�%*��f�Ƒ+�-�q��U����d6�r������q-7�g7]��fBj�A+6\/��.,��?E�9�*����U�W7�����ɽ-�#�5j��J�pWאT"WJ!��r6�b�g	�,K�G��9h9������v]
�ʹ�۲h�X���:�������0��Gܥ{cgm�6���`�b�^o���g]�K�֜/r�@<i���̻$Kxw��E"L���{nK��w!V*GR����ԗH���ы2i�;,�zt���J^?�H�vε+'�7��َ�d��U�����9/���a����۔���>��w,���~�U݆N�W2G��
;V؊�>� �W2*%��P��vY�G/��6$J���%�	B.�<��W�/{
�]L���	'?Xa8[x����@�:�������G�rqw��`��௟2�A���W���5��k��/8Gj��p{��J}l�����=3Y|�!�pko:@�x�#VU�r(�3�M�;��Q�4��u�,`�jg�`Q�ǃ�L�
=o&�*��M�/���ɳrԀ=_�W�	��[�I��&�f���ĥ��ͨ&3��?�T��3�r�D*sʔ�qi�d��>�=� bf@2vGs�����k���ip���~o(�L��ڊ�G���st�<�J��UZ#
߄-b�~�5h�!�C,}W�T�rl?��BT	r(���p(���W��Ҏ�R'H��d ��W�����_f��v��'�y8���j��m�<���'<�bN�,3��N�������^��X��Ɣ���T9߇��7 J�%�q�v�����~��O�{�T��[��tu6x�B�������8����2�-Z��bP���̨���o������m���F��m����6˽`��ʪ����#��P���k�ǚF����6��D�F+P.'���Ho�oD����F��1�S�kOxX`S'�Ք���;> ���|&�x]x����=�*m=�������g>/=<Ӆr]�F�_cbQ$4�_C�K��'��ٍ0ٰ���Y{�k5�i'.������ʾ����Z�((J=��aӄo��{���񼑭�99��a��e���^��\��*9�T
 .�-mjI��I\GңXkyD}z��ϱ���ڏ���.jC��߶���F�⇪�?6��`��9�$�jY�D�n��ݲ������l_���������-
�>4:3Q�ISL��]ǁ.��P�s�فy@�F������|��us�����}y� ~�ql�;W��Z�u�̕��{cڷ�5�ѥ+4mS�P6ju����`m���!A`��i/�:A�{��6=��Tխ_�sP[�"Lm�+����KW�F{î���S��%����9�g�oj��$ct������zs��y؉���B��� y�����57�}�Q�و
�:N��}�湉�[M�0`|��c��Qs���bOM�\��o[;�BE.��J�tt�x_�DP��E���'e�?�C�5}���!�Rѯ��aoA�Zr��d͋�1��Mn��1��c�|ڢm�)!�&���Ws�LW�f]���O�Ta�û� �, ��m>
�B.|_H�=�4�����Me���\�UQ�� #�2Eq�H�	�rNUF<�?��GP",5�_;3�1�^�0�U&����A���a�� ���\��d�m>u�~�"�_IS�z��X��z��:TZ>{�"#L¸�ߐO���#<�e2�M��Gnt:7q(�I�s���r���=\�:J^U��dD�v3��� ��ϊ$%�V/y�IY���P����_7�*�os^4���G^Ē�i�4��}��h��^���/ǽ��A<�/��E����V��l;�r�
'���hy7�IN(�C?%#��9P_�2h�|�zb����j<�T�-wz�(t��HQ$"~(���"G4�/������w����ej�e�|�B�mU4vݡ\k�Z�ҙ,G_ Z�A�����j���3;�@ES�e���"o���+� �h��^��Ph�Q��zG���O�E�/��(�� ѷn�3�_����ÒCp4/"Tx�e�^4!�Z��b�������\�b��W����P� 5��O���o�@�?A'��	K�= `w�2�`�H�!��Hݯ����"�5()�)m	-G#�;u�9��Jgݬr͛N��)�z=�={�s��_.��/��>����eЦ��>eT�������'F�f��:ktM:
���}�;'�>�E�K&2��T�9?�m�O�%�P�G����%*;m�B���.|�����9��64g�}?S4���� �$�2S�9B�P�m�h�s������P�v���Q�-�����h�hʲzM�/E:!��tU �<�����r5��>zB\�t�jƸu�o�>�ҽ�=���Sg�=��%��<J�Z�{����l�ơ�)�����/�+�= �FWǮ�H+�)��}����|��Vd��'ɥ�{� �o�$�b;���?��u�PGmt��:���ϴ|�E�뻙c��rKBt������wLfO�o:Wf��
ַ�c�GU4i�e���b���/�4�2KmJjms�9#����<!4r��Ùu5o#bQ�m���"�צoAk��"�S�aYf����ޭ�tm3�}˯�a���6��P����t.s�D$'�ϫ�^� '�l�S�D�n�v�L+�p؞��ɡ���`��W���
[�Ox���U��3u=�RY4�jb`�k����;N�Z���� Ǳ��P��!!�^cw��(�0�=K�������%���֢Z8/�j��^���qğܜ�Z��@�a\w�+Q���~1��6J�@4���2���ձ�<e��M���G,��Y���WPU��"	���$�i���~�fV%�O��K�6���2�r��H���w^�f�Z�,���6N��X����j�t��|���Y�П	Q�^��KZM�%Z�^^m�5��Gp��q��w5�d��&].�7�H	�88!܍u[[q|ly���~9�\�Ӡ�z� �W�W���_Zrm�!g�,���2W�&r'XgR�B�W�ɪk=��\gv|�����D]��x�ȷv��\�a�X_�f=�jO���b�"s�ATOqD����#���Hi��ήh��R�L(��͸�^x��ui����i�IZ�rp;�Z��+>���5��4��	_n��/��ϳﺬ5D�O�B�M=eI4�R�]�+GOWF�:<��]ր��mJ��A�|îRa�)��ݝ�P�����T�*�/���=N���4����l |\	�$fQwڔ���>r����)�@�UM�츽?��!��5�p��ܳ�6)�Z�V+�-P���f�h��3��Qg���P�h!�q1��E��I$�H�w�S���0+��i�7�p?U-�?��1�A���A��1���T`���?���:&�qO���L%��Z�F/�]y�Zr�	"��u����d����l�>�R���{�(Ay�y˄ȗ�%X��@�Z���j;�
KP��a�ݶ���q�R��-�� �;d4�4ش<�{�?oW@��ҧ��̀�~��� `k4��m�Iר� ��bs��P[�r��:\��s����A��l��xpP���5�csL�p�E��q������4�V�q�n�{��2��Aɰ�m�&���c6w������Y������`�%d�=�@��/껃o8��l��0(q���.���	�?[+[�l��&�k���
��p����(�it�����x��OѪ�*nJ�\�N��o(h�g+��;I|�����J�T}uǓ�4_{��z��P(*Ύ�Zo2�cP6�kM�f1���?:;��fP���] `���4��]���ZA�X��cg)�=j�]?���GV��D۱ P�<�6c"�)>\	"�����H���L���D�CU��{*�$:s�I3*�C¼�J+pʆgG�߅Q�_S6�V��@��`��I-��u)c���l�%-�q��#��^���H'W��tf�LCI�ܗ�2)��[���T�v!v�5���P6�$�<�;��М޷��H�|����p��`Z\)��tH<��|� �yH}R����*�p�,�G�6���H��]�ꫜ�w>�K^�ԓó_Tq;׶����em#@����9�}6�A8�4���N��@�T�p_����op�l������.8��/^5C���a}@���+2C���Cx:E�� 2.4����""��Rv��g�He��*�v�8sY�x�ʾ��GڵY��P��MA�/]�|��L�r��H���a�V;��� U!w�#J�ǧ.[�s��y[���,�A$HQԴ�9��,IK����WrΒ�P��Y�ݑK�@�`�\�y&�_�[Z�.o�� ��
��,�0 
m���I�^�gZXƧYM��u�}�ӿ2ޒC]D�f���jc
Gmz��k)X��x��Ѣ�E
q��=����u�<c (�ͫ��_�#~9mf,�+��挼	r�gL#4����e�A��6�<�hД����b\;
���lթ�n" ��+
>$a��(ǫG�mA���͂�5;���N�w�R(+5�B�@�G� |;�,�|}�����ݗ%8��+���ʨ�Nڈy!2� 4�{meM�L�*	���*6�N��6����Xv�Ԋ�qө�3�oXpu�����:3����:��c��)v�0�����z�8"1Q�a�Ar���������1��7�JDyS�w����� �`�/��g(���uHo^H���f��g�{��-
�� ����b �*kcc,�Y���j��C�����,�>T``8����ܤ8�Z<#yxA��s�W�\��P��ڝ�	{���� �����t�w���c	�̢��xhzȰ��h;���<�t�.���x��1k�d�@���G���M�m~j�a �ZF�xO6u�Hc��r�}��5xM�̻Q�`�葓U�L�F3���=�k�H n����u'�|4n`E�N�L�;�W�$j����#�/�	n�T{Չ	;�LIp���=��mc�	���J����{o
�;0�g�?:֭ޙi�F�l�����a������}���*��dZ�[�nr�▗Тϋa2�cFxo>n� �hV����������G��#{$սV��m|I�ߵGō:���֝�P��T&;b<��)��{����c:G$(�U!26���\�TaO!�;9G�p;�m��kk>��s���A��	�#�p��e��a��s��M��|]�e'�:�d���"mbs.�&$j�C�ª�@I��8X�^)[��z�1cՍ^�ў�n~	W�<���p٩��Kq\y_�'������m��ci)���T���A�.I4z��7�����h.e���%�L{��3���b�8�h������@g�,Ӑ��;�4���6��0��*M1d����l0����%Ǌ��{��7�K�i4_@ڝ���p��nP�M�?�z�:�V���fʤIa)��y�f�i��Z���A��	9FB��\�i}0��r�Mf����T�M�(�Vpr��e��qc���m�g,�j��d�*�S�
 2o/O�
V�D�O��h�ҟ�T=�<�p�f�d��[,�ԷMmr���	`Ȳ����� �Z���h��_���vi=��*A���(��\nA������\C⵨g3Iq�n�΋�vU��%�Ш|�ӣ�U0���w����q�0�6~2*a���9��r�c��N��ܷNp;�zǝq�\��B���'o)	(�y������K���}�E遒(~�~��_�g�0��I�&���R��1ub}8�_��	�ñ���&�e�܋�ι5�D2�-Ř��QV���3}S��7�k�UdU|�/��
�r7�:����ˏy��H�"X�Oڃp�6+�M�v����#p����[<)	 �,�5jФ\ǕL�pӛ��nT���A��Ք������Oi�������bNJ �5P���5�0�{�f���>�QC �2�xH�d ��	\���-Ƴ��(���. C������)��AV��_����N�U&9n�����FO�dV�)��9����� FԐ�ܲ�v<eeN�vIGZ�2������c@5��~��J��$��9Nt8`�R����6f@���>������s�Q��y����E�56��R�@��Q��$��$��:w��8��'����WC�a�v<VZ���7�\���&���Ly��R���"VrʂA�M6�z,��$�؁eb��lU�ߍ�I��!Q������gT�����+���O��4�n�x��̵�`���F��_2���E5�����D(p��ۮƢl0>��Ğ�
��̈12��I<^��f#3�Wն�:���?��{PhID_�֧5	����ʢkU@p>�G}�:
�v�9��x���grm�7��E�J�2-%yfmKH(�5?�a�
��o��B(�S*��W���B]����:���#2~��ҷ�S
H;��+֙�:5\B��c��Ũ��K�͵�lR�!����T��d�=�L?�<$�0~Yt�)rҩ�f�_��B���� �H���?�芫��[�m=���+�6a^`l��,{����_2���iY]�I�t��H؏�_��ұ��2[���f�]�;6���!���1�����v��o8�ܙ��;�Zse'��>X���jrOޒ@���gcE/��Q�oA.��'"�6?��豜K_���#�c1�ni��긯PpQ�+��v��Ӑs�_.�Mɠ�T�|��\�j!ɟ�x4�N��q��]���0#�(AǛM)�On�W�]5d�X�j�j4�M�/gZ-�|ĩ ����ZmBL�̵�6�|/�a$	F0Kt#O��5|�}L��*?�^Q�Uyqyi�]Ʉ3��"V����UZ�􀼘����6B{>���
6IR,�1��H|P?0wU�*������\�i���%��v(O��큵dD+>4�F�� V�bc�ْ�|��Ya�I8�T<����٘��Wǎ�1,g�5 �}�]+����Ր5�X�=��wX�;p��P%�����A�%��P��Z��Wo�e9����Jj68�c���cq�X��a��1�	4�� "��y E����ٱ�Q����r�zK�3��Y�k��i%<��n r@]D�!�E7��o��~E�G��L��}�EB%��t���B�9G����`�O�Wk�g����bl��o�e8���� �&v�ǖ�ƴ=�-q���ު��XֲKlF��Y��㣽~3��3{U>�&� ��5�z��-i�@��j�%�;̀�7�8�fC�o(j�˓L�'��U��Jϫ��J�z{̊�Xg���V7�߭�	]�M���>��r�V�	m�Qy6$�A+π&�S�d
��px�QeEwY�#��q��`O���~̊q-�菻������?|��� <���c2�����(��f�7ȴ��:�����L�������H���S��Lr�у$�I@���m�(�ɝ�FO��m� 
�U�4Y�f(G(��yh���Sn���~�g<N�R��$QZg��0�'�%��������>`�-��0ȳ:)�y���r(�u���������4����%Y�Vo���ʐ!8^sҡZi�����B�Z�DhYn�ʂ��A�Z�C���#SG�c
�>��{N޼����1�g�$;������;Qg�v������A��� �o6W�A�GF*PG1N��3���1\�Gf���_����K/LMc"��Y�
�W�$�j.Ҵ(o���n6p���@֧w��~�ҟ��V7�I[�y��фk�|�	��Eҫ�c�f�^F���Ͱ�dO�OuA�߆�8.�~mgS|
I���%~>%bz�.��]:)�#�o�2ξ�ɖ�����Qv��D�9{����Vn]������Icv� ����x�fv��S��V=�����mN�qo�~�)�x�[���g�iT�WWުʋ�!6�,c?�O��*2qz�W��y�9��r��Mx���DP[�*5\3\hw����`2M����C}u��)3��vV��x���3�
�0������x�$�j?n�I ?XI�r�n�'EKs��H�e���G ��丄x�e"f-we�8.�����mCvT
U�91P��)���i݌�R=O�h����>����b�9�*�2�ȶK/NI���S��b��X$��gh�xt�WL<�2�Dڽ����oSMS/��C����@�D�@���.� ���#`P������pݾ��qJ�w�Q50�c{ґ���y�6((�@u�@C#�[ ���-��Y�N�u������D^By���3�5k+��l�L�v���fW��4e�g�+��[����*K+����2��z*k�hٚ��k.�MZ�NG�ҳ J�Z�c_�R��W*��0e�CWb,V��18a�+��lӲ`���
�.�ǎѠ�ﵱF�:,�!su�eRVjډ7e`����R�_Sݡ!�sa��DV-��l�HyѨ�?�5�M"O�ȝ9��@-�Y���Q��n���-�O�<�'�����q���	���[5
h��@Dwtv�6Jg�D�Z�����bdKd'���^͘��5�U�`�(B�Լ��;��ۡ[k�dO��ͦ$��;�%	:.U	�[ǄB��zp�y��m|D~�B���E\q.���+�;�I�e3��W3�2�o*�7�=�C�l�=�c	�Q���!N�3f����d�� 솄2.�	m�A�� ��M�����G�{�c���r���J������yt����N��G�O�0�+R�y|r*���O&F�!�V�[0� �W��_ʍ,I��y���|�6�����k�,8M�T��&��1�a*|�,�j-����ᅓ�G1��gۧC�1V�������V4����=�̩)v����o�IM�l_5��
2V+��t�-3^�����)�����J�1�	��A��m�8��G)�-g�}������n|�� ���ʾ�.�2ӡD�.�Tq�{�����tQ �R�՘Q���gX������j㫰��ڿ+�D�x��I����(��:7
f�8^���}@������g�$"w��	�bS��]�ű� A�Q�R���&�w�PXR0dF���M�oͿفٿي�N[4�b�����++�&0�����Y6��Bޣ��?`�6{�LЋ6cbN�HtsN��eU2�<}���r"a^UL��0��KႈP7��&o{�U�������,ϧ<�p��\M�2"���>�gQ�~�r����jF�tl+��,��}U��0��53$�V�����iS�<;�����]%
�H��&�׏�9�l����6P.�Hۂ��U��D-<�bM����I昵���%��j�Zg�,*�ϬG�(�vs���}���	e�S��N6K�@`=r�0�:�3�ۦ1���"�S�&�"���*�S��[��Rݪ�U��$՜	����p����,v��� BC���OS�;P��M�b�<���
{;�k��=����β�ƛ��)C8[�.p��н�\����f�^O0�4B����kv�v�n�#��1��p���z���I��W�.\�V��@�����V��;��4y)����V���g��]����.��=#4I�Y��;�����0Oi�h�܆�9�7a�B�o��d�v &��"W���I�R3v�4����}�+��^���f���_��\ψ��W�S"��_�R�V�|����ݭd��X�a���������t:�j�BV��2��əV�>�x���j�D�P�eA��E�9�@Z�N��-��Z�<���{ԇr��kO]�|�"��}V�M�65B�� �OV�s]`�����8Zʭq���w��O;�T����ކ�A�P��� t�Y�#^wQg{�d�l�
�^��פ��/+)s��z�i������K3�*GT*r�_�#.֩\������e_�y�a����gb���5�� �`n��������/��x1c^��6�%�i�@b��
H��KFIq��3Q�r6d@3������������C�q1Ͻ�NH����J4��,���J�s�5���d*�Y,
�%mS"�c^}GU�Z���}.R��~��?D�\y�j(7���,����x�w�l�X9�}�����t��[L1H(�� ��tGH ��G��N��-��)�t��C�x�K�59#x��P��B�S�U�"��w��l�;{=5/��{��
�e�ze6<��Y��p�-ZE�"|�
�.�ЭLv�jeb$'@���t-2;V}Dѩk��Z�;����c�ڿ/`���.���q�6���j�Y��b��J>_4"�1�� �F�s���n���p���ǮmǨ�� 	�J�6�n��3�x��+%i5]9&��p����.�#}�T7R�+��[7D��S���' x	.kBTZ���^e9�PǒN�[��ݬ��+w��3�Ĕ�j�9��W+2i��K`�Mu� ��m�r������I �d���Ǐ|J��v#��fD$I��Ǫ7(�3,DI�i�lQ� �X�nw��YRP��9-�d��:���wM�;^K�^���@g�S�D�EX��:I�#�
�
Nbwܥ�bH���4�{V��F�2`��C�B�{��j��ߪ5uϱ3_,䆜�7��'�;���Z��������W�D
�fԠ�IEj�gL�V��@��g��d���E}��:�A�b�El~
cރ0u�͹��t�47��C�̉}�2[�E�;�O��F�����Iq�ZZE�;XL�W��Db~Kn��	�ĥ\ú5�C�*��0�����>e�#�|������	�?ȟ��T*z&c��>t����gK��P�_��R�@�B_��9��q�B�Q�	0F���5��E?q�=ӓ��kD�^t��Y��0�r��,G�6�j/���㒹�z�ҷ��WJ�<_І�~��5.�r��V�fݰ��T{mb�VԊ1��$�s�g1ߞ
�}�!��*gw�4�Øm�V��`� M���%*�S�k�7�ą�EI�pU��ӭTO�NC�%C x9�/���Ē��)���x��[�oJN@[��=6��t�;�� B���*��M�۳w�D�|��H�_��[�M�$�|h55��U���͂�*�R�@���z�6���P��T@�@��	ȉ�<�����d��x��ƘùOe\�j��g���1b�iO��ϫ�T��g��Ka����ց:ݛ�/҇��)�pJK��z�m�f�r��G��{�6OA���K6��� �}G>َ>�'@2�g\n8aA>�sU[A�q���:\�+��%�"�!�O���r��h׭ۂ#n��V��v6�� �~��������:��,�c�����A�Ǔ�8?����̤�Dj4st�� Vȣ��i=����7B.�}��Y�0�j��*si'd�<�9ؼEM�y0N� yL�/ֈ���[���k*8RA�.{���D��T��f��eo[���=�+��N�,}:B�N�y^���玥�<�4��
�,�nAXQ2<DE��A��?��+��u�� ��>N�TA�T���!�N��`�{Bb�ri����xmn�nm>&��"�yt�h�^�#l;bz��t���-7�\K+�2���'�e�F����'g������J��+C����_�X_��cl�!Y.ŉ�؆?�J��{�T��d�:AX=���(P8R_Ws��'0���] ���h!i}���q�Y��z�<$�)d!�Kr�kY��z�
�/���强�oȨ�^��,h|1�K��S��7���Fܺ���oW2.S��_��ѼRZq��<C�3v#�.�����Y�`*J�����.�6B��ˤ��a������8XM+��I����ǌ���*,?8�_+ٴIQ�P��넨Ǜꆷ�c��-:�h��S��J(�O����5��v���n+��. ��Y�<C6�1 ��|�ڄ�4�@�%q��������2��Bw�b&�*J&�Ɵ#��vԒ)U9�l�!Zg��p��K����n<w�
>��&��Q���ndk�&���>K+{$��O��Y>ҥ�Zu=Se9�m��b.�@��V�/��T(b��ȓ�N�Ʉ��#�a��F�_3�9���*( J�;��)q�:����
��#A.����cm�ax�%����T7G���P��aC�>jO���T�Se�J��P��Ll��Ez�ob�yOr6 �k����+�M��c��?4���Bvf=�͂J�ᙃ� ;T���0�Ϭ�+��x�iZ^
|�T�}� ��>�H�Dk�D�tO{c6^��-r����j]~��I>2v	��)���v ��tP���25	��\�} �i�O��f5eHĎ�b�g��i0]GL'����X�[����s�J�3||&��GH�5O��d]QNJδ�!�y�^^�'�i���?�X�p�D�fqT`H�'xJ��,?!��۲+(.P\�;�;Tݻ��m���=q~�1_9֧��zL��'����չ��j���x��:�'sf�L4��ş��*�E���?0x�'F����=b��
G��R��[�g\G�QiC��syk<�bǛQCE��d�]n�[l#��n�k�
Ը{7�ѽ����gRB�!p�Rr  [x����ʷ��W���_����sV��b�d���Zr@.�et�\l�o�jz�׃"�a.
S�p�a�����P�(�b���.�?�'�6�WC�dH⃞�T�mKDb�?�%����~�� =ﶪ	/���[Yn��ct�h��YDS��b�j�-�c V,��/7�����f*��_�=z���c��؞y�Ek��p���<3��x�!a2k��]hѤl�~ũ�J��܀��"|�6I�VE�,��2�}jW���>�DR�`ƼQ��e'����R.j���{���)8�5�����%�������md�BOAmύ���������������eo�>E�:z&���`�v����N[9�����#�ـ�1������Fkw3���w���	ʘ���3��4���\ؙ��\�2иw��з��<���#Xr檔1� n���*ܖ�A{ i}��>��f���y�^�6A+s��&n#�+�˔�o��:�`������8 ���%��i�5�/G��W�_*g�L6=�pY�33K�@��M���j�\����b]�(5ca���˝r~�9�D0s1�j�Ԁ�Y���� X��K���=hm�l��K2�F42�h�!��H򷏐m�\��X�0�܌谥���D%z]T��Ȓ������8�p�(�s����@8�N�IS�wM� ͎Kr%!@c>^�r�L���;@ �Q�U�x�l�`�P9�w4�5�܉�ٚ�����,fY�w5����A�Sx�\?)K�gau{S�@�M��"Ԥ� �L�ӈ7)q�c�.	Ļ�xkj�a�_�?R.y��Y�p�Mf�]-m���u��i��ݍ��&	�,�V!�ҧe�ێ!V��B�Y��&��ܗ�*�݀�W{�վ��%�R��wQUG!���b��f������A������/���V	_@C
[�� Y%%f9l2���|�XGSW�2������ϕ5{����o��{�ɀ��s�=��S��I�/�{f/Ɣ��gJH�?Kqy(��	�׼}ZwVn87�h����h�u��Χ�m�����Reܾ��ga�!��W��H~0G��蛕y����|Ά�����O���@�o��:���gᓤ�T�ؠ��н�m^�yR����ͯ��=`�#�i+#5�����s9СH��gR�g��!�-[��L�?ڸ�c@��9)� �,c�B��O�ғ�[�����o�U��8.�tҕݺ��k�nP�]��q�u{k��k�L�<H��Ps�E�t��wn%��4A6�?��0�J�
L��������||�8��s��zf����[���a�x��io'"��~����B(ȗl}6AQ�wW�|R���6�����ہABXd�h��T��ِ��HP�^��%]D/��thmT���ѧ
#l#�
\J���	���.��R�9zq�ྷ$�̉��$bԵ� �,����0t�2#_�t�G������A�����ןsl�woDꞫ��G���.�����;5!��4��y8W�-+i�3�����㝙�����4sV*����#�=
��CH'�1�^x�oY5���Є*H7�cՕ�P��ƪԦ��ǐ535���|�Cr��tU���ʭB���z�fv�Z�����ia/\��m��s�+���tx�.M��e�S���-?�����I����#��h�ٟ���cPC�����M��kS�p��&v��
�u�����2�E�	���Sُ�\��x|�/5c��]��t�Vcj�
�	):U���U�̑�W5�+�2��B�2���̡��:bz��1*��/��H����K�q�?v~�p�=���N�� ��c??YQ��{H��2:{*�Z)�I���t%�0�Z8Cc]�гv3��k����'y�?�y�����X\HAOz���'ݝ������<�4��"�!xK�"��_B[dH4'����L'b�ⱶ�)�M���?)�4��r?[�@"�së���OX�k@fAy:�����?�^(E
2!�kF��(N-����Ə�r��S�*��3�\�//�l�2���ĺϤ�ݱ�ɳ��^S&I��c�a�Lǀ��Bl��Ht�2\U��].|�k�_�DC #�<�&]����
�|�`87n�����l�_"��Fu�s����2������*���L��A@*�Gt�F�V���W�ۖ��S����a#Pf�?!�8�p�4����Z����\�
�o�h
��!��
����v���<�r;���B�0R��{�����3Hn����5�y�5�S���W� ��w7��㺎�ͷ�>�V��� Z`�zHC{p���#xj��c'�P���1�Xʿ�7��^aB˓��h���vJC�4g|$��Cp��N|S{�+g�H$[Y^��`�n ~��(�����Й�-(��
��������t�ī�����w��?Q>�l'���Rk�RK���L�5j�y���0E����d�o�5q�f�D��-0�*��)E�zd��y�s�>���7��	�\+��͸���"*�o,v��4R^/��E���{���?1n�UI���\� oCmy�'�N��!U��dJ?�@O��h��Ӕ�����H�ᦣ�K�5�RBiU�C+�g1��=�>�ƣt~'������O�f�������\���yc	�S3�tXɛ=��2�ؼZ���(�]2�ݒZ��Wx(��ɦ��ۨ��pfy�?E����`{q��/l8 �Q�CC�+�\�Y�r+�7��)Ԧ0o�Ld�\���D-�l>wB��j�e��'d&����PC���N�,P�ލ�x�&�OS(Q[�������P��ԖF�}Q[�<��_�W��W�L<9�sH��{	�nZ5�{���&R��b�����p�ׯ֚F��C�#|�>`���#^[?S�U\�_�wt��E<��S��ܷC7��#c�߶I�T�����P� ����/��Mt֝�x�!�KX$§V>�#��Oщ��v 1Y�b��k��RZ̭R܃��=��nt��-71�uO#��%9wxg9cfȧa�>��o��Ɐ͒Hw����/>�O-X.�U]�6���c�>X������[��?�~��[{M\�����W�&5|�ZS>�m�����Xe-n`���2\�9�e,ɠI����)ϭ�A��*~��q�T��Fg� �sjD����ˬ�*�2�����*3vh�'�Q��T�U�䗙�׭,F��VI�!L�k"n���Z���bcRҘ�f�JA��A#_���ڿ S�T�J�@��ue�L%cu�4ᡧ�S������1����R�k�U����Af�x]��O�r����Z,�&rx��7���D��� �6Z�sA��%WHy���f��c<�a#�y��z��J<HE��$�SHf!΀Ѫ޲���䛋��D�q�����  ]�V�Y9S2��� ���\��λR�ۨ#,2u�p���$F��*#��|�f��Z��Vm;(�����x�� @.���w�ǓOǵ�����#p^�u����}R�D��2�y@��`��bQD��W��P.	{�*'�,j�ĉ�����F�O��*�qo�7YWe' :d]�jS��L��g�x���O�n����m*QU[�U��+/�X2�x�vp�5-�ʺՇZ=�ζ�Y�dp���)��Y��wXh�ᲆwV1��zk��O>����vQN{��C�%���ꄠ.�J�*ʏXl,��o���,*���0:��
-�`�y�Z��a� �0S�{����z�"�$�k���&�2+\`"<J5҅�I�2&;��娑xD�T6\��5[L�G:�'ƳD�°J�yԏ�GLkS;z�_�["�
���=�
�只ɩW��* �c��&�5u}�S)��ک�@k���o�S��vX�2��t�eg�ژ�H����x��G��:)M�tbV6S�d6� �`���>��]su&A�Di�a��9�:͘u���Ex�>ITt����i���.��A�LϘ�/{��K��? i}����#>�C���d�)1�d��+��������NL��eT���{fQ�R���spZ+O���|Z�K�l�`��8��9���tN��@�� =�U��"�<R�*��Z�Zu����kD\�̒k��s�K�jI�i��Z�����]c��'���=�"�U�f�ݧ�#�`���G�_�#:�+�Q€��ޑm�K*L��C}5��k��C�~��/�%<�>�������B�X��!�J��XO4z� ��L�J���#XtH,�K6|�* �>����e��`dos�����0[.L3`��40�B�W�P��?l�3Q� �.�O@�zG�u�_c�+(���7ߴ��,h)h�n���-�mU�A�Az����i��Oj〯�1�7��9-���0�#X0v$���J��&߂�e?3w�p`��Rǌ����C:u��m�!u�� ���f����h�L4�`��Aǂ�g}qr�Ĺ�f[�'�
��Zuf1�wJ��K�.�ه��{�T��e_f�K��H�&����5�؝��w�>�+o��NK�̯v8�]��`~���j��	��<+ݐLǣ[f��F����
����4���
�
L�,.%��;b�=�;g{J��d?�$�jѿ$�w�G���oӑ��DZ`�.tLu ?bUgЫ��T�Jp�z��+��mv�uc�Tc�֟xG��i%����~��o4&���6�fVr2��c�DcJ�.��gէ��ғsN����5��l�Nt�l��N�m�6��w�!J��6�=v�.���Pi��Z5C8Q�����ې2�m���#�<�0u� ɡV�D2�� ���cVh��.��=]���};��u��f	��x5}l���]��O'r?D�Ll����N15�J����K��G�%�?��������n��w�K|/�����{�M�?��7F u.���z�����ܫ�	������i���d��ي��O,ż���Vo�k�d!�o�fjg4��;�yQ�"���
�F�~��8/���j��Ù��[բ��i4?�ěɝ^��pCpNiNR����/[���[�Eea�)
+`�h%Ƿ�����ΰ�#֟���m7_�����.�0�R�l��ɽʉZ2�L ���B7�E�"���f=���bUW����:�q}R_�%�g����<�}K�<�d"m&<>�Zn�@vj�7,uW���pB���9��q6B�S���3�z�$֨����9���t�%��bD0m�)KN��BZ�j��;�S�ɔ_Z�:��U��-�r���8��&Y�����S����B~M�K����C����֩H;Ӳԫ�Mo�;��`�R��js�p��^��"��� ��ɞ%�|�O}�����YV���/�x��9�Ș�V���j&�˅�6T�J+���D�U<sP�n�`!|��z&_��-m�xT`���Qh:c�����\Ҹ���E�:��X��O��aq�P�,�<Td��䜘aԥ~���{����n��|�j9��B�2��`�{�S�/��el��2y)�G�~��ѓ��\�y^�htO�oƦ�ۋV�F�U�k<_��k�^[�������)�Z[�.���$�! *]Q�����M�c�9������'�=��p��`w�v+���X��Ume���������,�G[7�XE����͌Rok�玖SZ���5O���+�: ]y�\Ց��i�5�$̦uxGO1��#R-3�Ƨ$�#4;ґ��t�[�u�"#�>��]�O�"�j� $��w���Z���8��dI�B�y�O�dF�Z:�y�E&y��u�bp�d	#�J�1��UtgA�Y| '���\Q�:p.�!��
U	���k]��Ed�v��+�/ý(ٓ�z�� x'� ���_��4��H!�8|Qs�F;ϽQ�M���KZ�����:������Y�D~��h�PV{%;��w�&�C�s�<bϞ}�wX����f��,C�O����|�ئ/�t�w��� ;�V���i�e��TY���]����;��sւe��Mc����U[Vf\��P0�W*
��#�-+1�
K0&U�oz\�_tW}$����d@�_�M��ms�㞶�؍�m���V����+l�N<�<��<՟-����b�ٱq�G�Q3�ea���.ɒ3%E����K>*MfU��v�q	��7xB�O;MPE$�����h�R��wIl,7+�;�bگw7��`����b�:�c$�7m;� [g.BeZ(�������w�_��Չ«�l7��E�MM|������L�$�f�N����k�D�]���{<��'�	ˠJ�������E	g	�bcE����>3i^�O�Ai;��N��s�+���@ם�#�ovİi�{m���H5_K�����^}���[�у���K�d��γK^�ϺWH`kj��ۭ��|���Ut_a�\�F� ���&�V/AQ­��%�t�� ��Zn��8�mi!�+^=�=�����B���h������B0y:��ȽeU�j��Q�jf �Ɉ�H�"�Z�Hm
�����������"���C.v�l3;�$��Vf�U�b0�̠�$݄};�]`���t^�_չ=v�cf��t���L�1��M�ة5\�(��a��䖗FR�ϦMTDc���i�i���A6"[��K����/rV�p�^�ӽoB�׶ }t@��f�*�wb&�4ͨ��9��g���pOZ7y"f�"�Pb��I#���
��/��/)?i�E���P1U���L=ְ� �f�UI]s�[��̢���*���Վb�r�:�J[f�Z�\��h��+�N��(�
)ҹ��-S2���ҶH.p�6�͢�ԠH �x�	n=,�eC�K�ݨѮc��&%���h
���8�w���t�$'GI��Y99������ ce���S���X� [�{�<!����;=�V\r�t>��.����n��Rak���@�^���M�����HB����í)�ݽ!QhȠ��K�y3T�ԡ��g���A�<���υ��A�!Q���G>3{�i�g'�a�D���2��4�����^,C �)���^�a��D%� $�5�؃��&�_'1Y�=���s{ M�x+hQ�.kx�I�(�}�)��ؐU�h� ��l�٘����yL=?5�i������
D�f��h���X��)�u
Xu�0&�k��7�Ud�� ���Nx�}̭�^�r}�"���1U�B��c�6�>�"`y7�)��є���nԩ������f�@c�}hIs����/L{D�����L�_[�8��T�O)���meWzl����e�����a9���a�%�����6�Á��,�"Ñ��+{܀{����`�}m�&���|�s.��%k{9U�a\�8�+_M�u��YG�#��ɏݤ�G�5���?�Gu�|�	.
����Lk�����Z�B�	���p!��V��M���6�J^C���(
�A��u�¶����m]��S��e��	볽q꤄Е�p�͂O4�%FU�i1����L�9�W�_x��*�x�}�(V"�ք��5 Q*�RP8��m�P,7fL �f����c����8h�)�G�F��kBq�<D���{�^�EzXh��{Ȓ	�]�;Ø�b�b4�O�X��ex]��<ηEj�%�Se�v�s4y {�T�	�_E������G������ե"��`lDb�E��	˪�^A��Ż���L�j�����/ƿ �
��##����XMT-
�V�'�Tz>�z��_�ݼH��2��pp(�K�"[@~/�<����]��\+�}��ڏG�ү	�ԍ��=�p .o�>M`� �Tٞi�-�
���Ԝ *��LI,2_���R��>4gL���r��(��	R6!0�^-�6H]�0�^P+Z`��;T���_�<�b�.�k�>u�I$π�e$;�Q[
��?E����zP�発O��kwA��"oE�?��p�h/X	��MH�h[�8�:#�������6(�S� �����Z����dG�h��
�%���~f꽢�aw��6g?//h���i�; �ض9���G#��eoJ��,�KO֢�o$pnI�(9��܎��9�"�*ǘ���VV%]_���O��݃*����?n�.)���	��^�b^��v��,�`o\�OA�8�wJ��
��"�`R]v�+�8��땸:�D�����#�4fr�;+/��{��}�ZWȉd��pm`t�
��|y �0�zon�]bة$z�ܗ,��b���7������B�c�]QR���J�z��(��A��'�b��0�$'�����A4Ͷ�p[  g�+	�S�R�6V�ϱ%��Κ�L~Շ�=�����z��ɣP�汦�ı�XJ��q���s!�b��*,
KS��v��9�$jh��~�r��T5�9�q�"�$q��1���WB�Zٟ:�(� �,�1�~�"f���"&�k�G%�m��"0� Ksuǜ�w{�>��Nw�p��RW�����:5C��t҅_�a!ι,W�j�\��,�+l���s���i�i;�Irh*�O�_ߕ"x�
Ru{�a]� rZ��%0�ΆZ�l�d��J(l�X~�k(��3�Q�_�L>�)X��l��������c�6k�m(7��h|
.l٧:��5?0QE]ɳY@N�<K�镧l����+0mW���۸�\j�z�>4�8;C�I\�^�����4*Z���۪�mD L:'�_��FI5=Y� |Ý��I$�T_l�7Om��!�i9�v�ja�� lJZ�*�#���l���/���V�'8r�����A�!�����n��ø�%�1��+)����)�U��v��	�"J�����d�V.���gP\��bk��)r�����К�jYu|T�<B������Tڥ�T����k����2�&Nǿ� �6��|ZY�5�:L�Е��]�N|Ή�$�Y�(~cA)�kxI��rY�sg$�
�w>s)[O�p����Yk��� �G���g`R�� `X���	u�@'�b7�2�t����a����&f�d)���A��8�7�iT=�!�f������f�$(2l���~t��3���M���O��#:��2�l6&K;��.+ފ�_7�J� �)���-A%�3v
|����@R��/Tb4���2bTp�%a�����L���z���$)'����k�����]���t�5��g���[R�㿦%�ؗ>"�V6OB�z}Z�:�2�i���p��?hl3^�OOʦ�M�op�\�����v;�z���'�P:��[+���yQ_�^D=c�uh@�/���+#������6l�� sL�F�.^��JX�b� ;/�W��\|t�:l%'Vҷa���
��qCm۴xA��b�C/��P&*I�h������B�������2����D9pr��3���N�Շ�,��%޿Y��(q�F3i�p�����zV���1L�-�f�9GV"YV����q&?5�f�����࿚o�A�O ��??�w��TS�S�B3���O��>�'M�s@M�{��1s���O�7�ށ27�h��4�$�Jj�v�>/d��;@�蕭��l�D˪���LI��1ұ�w�	�%�!�),�M�im�[H\�z����:�r~Q���"T�6����-����z�f��Ĉ��%��&L�t�j���[���! ��T�qPݜ+�}�����ıR'�t�Ss]��q$G
��!k~��㓾�y�xV/y.H ��
���� ���Ŝ�XU�~���Z�*���#^�W�������(�X�	�.B<y�20��z�J�+���v��0r���v�;�5c�5J[ͭ�HJ��:Z�ޤ7]U�����"~klF0w%PF��,З��S2��tو�;�J���Vo{��~��%�,�a1��f�Tl�i/cwk|.Rb[�,��j�9M���'^����+�Ա�nRP�Jo16iY�p\!S�|�#;H�����A:5C _ԇ�.�Ϙ� c7� U2&7eۂci�x��8(LZǚ�$���b��ɉo`��eQ		q�8\�Y����,+M����x=),�o(�AH:��,D�7�R7��8S>���%�,y�j�[&�O =j���B�߹HќC�!S�\f�-�"P�V��OϷ��~��}��]�M��EȂT�`����C�n�3PQ�p�E�Z"�]�O�0�8��	1�������h�b�,�K���-�Jw�%8Α,-�W��,����s��@�xP��2���4���;-(��i�x+a�ڃ$��L��Q��� ��w0h��)��hq����(=w/�+[0��+��_�#e:�=���i��5JY���.-���>�3�݄St�G�6؈v�۹�J\��A�Z�b2d���e�]1M�$ZX�v|�&U*��e���3]5I}�˱Cb�(y�&���d�Q9_:�m� �M�	
�Udq"��q�5i�0\.�;�l�T�O1��0;��]_�_9�����Oa!$��h��ކ����,L��E胠\���Ez��0�Q�l�rL�Hӫ3C4����B��ip:'Y��������(f��*&����	ħ���}e�KC����krй���3nD�ElT:��F󹨇�bN�(=�&o=�(����&'�A�@�U)yWG��B�v�=Q8���!z۳'x�����/)�e���z�~~/���L'�Ԯ�<J/�t'�̋��se1�����w��c��c�� �*���W;;���ܽ�ر���iL�J�n=L������^�~��s���M�e.���KU�d����%�^m���\s�g_ܴ-��^
�r�2�yܑ.y�t%�op9#��@ ��3-�Gh����e�NC��6Y[ihF.}�os?M%n��BP�k;��3Ԑ�MNG�Ҁ<I��cD���Iw�gS܀� �o�k���5P�aFN��?#e��+�Ү�D��ŴK�r����Jɤ�7�H����^�5	�Z�A]%�H���b�����D��'��虺(l�2�ڑZ�;EV-~^�C{�a�c4�}?X���Ʈh��h����[�t�M��� �@4Ce,�s��ko����ݬ��KL����V ���g@äIoǃz� ��[ �g�8�$*���3w��t���~L�E�x��{�3<_�]���f�G�	�y���0�}������AP�`�3�����Z*����d���Mn�$�1��>�P��f����H]�f6�2�.-,��Baa����j;4�,��Ĝw�t{B��ɢ�Y69N�;�!�Yrk�%��1���n�v��|�I�ڻ:��Vz������~ژ�r�c��'�"̓i��(n(�,?"�D�"��J�!Ϭ+��	������/���Ȉ{D"2n�6��𖶕a�f��k��I�H�W���㛨��gq�+Q蒔��	Ú�����Kў�~��BiUH�������xs�uc�5|��F�dp(�v��S�S����Kl:q��3W��y�x���%S��@��E��)p���m.���Z6v��:)|?�����f��cs_���@ ~/�s^��J�g��w��<s�k:̬�?^������M�K���b �v�I�KZ�+�z�}_�wV�	��A�����3_����Pt^�i���x�1�e-ym�aܝ�ɿ�"2�Z���S>�h���w,*�%Z����zo�4�Z������L���68>Б��\�&�17�7�ݲLDOӉ�ȵBDm%� ����� |&)��
�8\iH9��{�8
�� h%I�.��~��u�������0{�𚹃�܏�m梛|�P�g�=s�n�U��#��%^cIg1�D���G�g�C�w�=��2;�8�Kmz1E��!~G��%e3}�Ns�!"q�#� �Z*u�6-����S�Ii kJ�X)���^�D'��-��)�w�?,�5C�6���wΖ>�_�_�
�^�c&�P7�{�^k竧���rIY�yF���_�.����%$��Lc��;j�Mr��.���j&u�f�1ߣW�"�L�&9�
{�*H�a�~�jy��zӖb��z���rOY*Q��ɹ��O�8��n�L��ݏ���li!sl��������7�t{tO�[���1��M'
��,� ���ػPX�^�2Y�|����L�l<���ا�_-�^�b�;�ҿ[��>x�0e�z�gs����2� �����K�g##+�l��C��+�z;�9�*����ډ���S���"fVan�J;�D"O��i�z1ν�(��vs�%U�y��&��8�mw����=�B$����`#� pg��^�H2��9��Qj^b�3�X�-�Ef�b<쎩�����≖��zVs�3���LH�孿��}%�� Lss�e�!�.���t^"�Q����?_Jc}������*��w*�=(��fO�p�9�p�Ա�A�Ş����G�FP�Ь%r)���Cir(󥜬3�%�f��9���󄑬l�T;�ޔ�D傲�R�n5YXu����UjS����J�`�`�J�Z�5C�6���ŝ7����)�zDA5V�v�ܯ`�$1�7��~%4�`�b7����� A�kh�D �BK$��J�\��i���-��@^�B��+�fj[[?�� �F�[�+C<��"�O�P�4�TTop6<i�g�ְ�:����rOT��Ŗ8B]� wȝ�Vf°Y<	Wx^�cL���߰fM�  ��Μ�*{�����w$9��_�G�Z�����B��Uvs�(��f��!��Í��5R��@�b���M>] �52�#�x�`�La@flɃ�;�P)���W�2D�����͒>�\�g����A����D��|��_d5稠3��I�_��9����*���x�HbH��U[[���&��2�>�x'�aT��BޭM�����V�KIZV��/�9k�"�����CZпFV�����;T�K[�W�nV� SuB@Y[L�`�������~(�� ��R��ɐ��w2,���۲�]7���X�5��A���L$W��z*�yQ��}�S��8�M�pyw�f��F"�ZMsL�\��&D���R�Lx2Ed%,��5�/�$X�i��Q�R��K�*�Qma<�#SD����iXdp�4��e��D��3��7����&�q2��+�7b���_7�323��؍�a*���֌ةղ䃚��v�ʬ� T�F<u�@�[�|X0�	GY?��e��O�o�osj*�#�ߞ~%m���%��ҐL�[�on��Gu�>\P`��8�Ya�<�
n���:Y9�Y�ƞW��3�w6�5�r��i;��[*54�V����!ښ���G�&�hp#��5�����s�>/N&���l��d��P�nTR���6	��#��8�v�����:�
V�8���)*�����yk���~�6y��k�RU�fKQL���"JJ�����!#��5XC���%���ߊ��������vU]��.��pn�n{����(b����~�9t���x�;R���md 5-������݀"��y�;:(�=^Q�q��1bd�;N5�BU[J��M��4>�\�؂��)�J�y5���g ��3ĕV�����=|R��BDo��w�r���eEZ8��KR�T��ۉ�J~�F�i��+�_����b%��b��{��ٌ�դPYB��j}'�����A2ي���b�<G�fKk.�<���$R�z� ��4����j>.xwQ���p{O"@�I����J����rY\���vx����q}�����b��Y2�d ���n�L���R<���m�V��{��J$�j�=k��٤�9$��d54IҳC��E���J�/�`f4ʻ���c����V��IF�ᡗpS��b�Q�f|�{G[4�(�_�}�����>��IՔ64Q8�ާ ���K��x�=_�KnN�^=2^#�n�T�"�Ω��\�6�|��Y�yA�$��[tS�m<.�F�h�'Xt�$,G|=��:�Eg�}�EH"j Z��S���r(͛�Wj��Ø��5�,�(��EQi���_��d��l�|�
V�R$qޅ�Pf�ꄶ���_���f�{�yq�M{L|�Ty�t��)b�(�'C�;Z׾L(vT��'+Χ�{�?�pCň�jw�V��K��4h�kh�&�T���'�ڪӢlD�Rs���d�+���*CY�%)*�mi!�_�m�󳞯�P�ɯ�}��3�w>�XI	�ҿX��T؆�K��u�cWU;0��%�3�^�N��aֲ֍��4��}��n��V����S�~d��������+�{�����������,V�i�ۓ2�_��
���觥`=��#�ծL����E��6���NV���5[�]/N�T�n�����P��Lj���A1|gJ<g�h�$���q��q/�?�A� �Vw緉F=�S�ϪU�;i�o�v}jҙ��K���؈�T38���`]��t��<���,���zT�7`��~�t�P�t1�&
x�A l$.�U|�U(��4_���]*!=�tU�� ׮�3���umP�Q&Uz�$�v�K�����t
�����H�o6TЌ�&Ѳ�d�!z/:|�=�
�l('��sy cK�����c�i�p�̪���Y��s� !/�y	����o9��P:��AG	���C>൦j	�
�T�憐����PR�c�D�34���0-�����Z���*��_�Ѱ�Մ�β���]'F�h�k��k�`sMC�Rvѩ���ӄ�eg�5������g
�J/J�ee7Y�e��|��-K��䴵昐:�C�z�o�+�ۓ��^&����0A�ԩ�Os_.F1��v��>�K^�
�<�`s�n�g�����=s����3�UVf�\�w�?j	+��CT��Uƪ��V�l$0g^��!�\Gz<�#�MZ�]�5�gr_��MB�w�&���h�4��d���6��?t�L�*�߈g_��HJ�[&���"��N5�6��F p|Cb�5$�L5�θ���R�S1��m�$1+���i>}��n}�G��;Z�bY��xy��q�~�O���gE��F�����ߛR' �����N�щ�d��]���F%3u6�R��?
ö����\+t|���T��J�8m$f��q�A�eu.X�Q�W;zn�������=㚗(�'�+�w۴�1�H_rU�:�ճs�h.�PC�	����WF���)MtP�Y^>]4?�:�C�1��Yi��<�i( �|9 Rx�Qf��-���3ʷ�Jl����i�]�'{�n�#�g#��K�sG2@�9��}���HF�l{H��[L~5����Be@�&g��_b������*��f\|�%c6�HS5BvWT��q�&*#���@qU�������3j��$R�w#l�.F0��K�m@ka��v	��Rǘwϫ읙}g�ǿ3%|��*�����4����q��c��^�L��\z��N�q�8/ó�#y�Uvc�+Keh+#��,)��S��aqM���V�������R�I
uA��c�_mǴ`�t����ͯ��>�B����@C�ˡѕ^��s�?����EU�:�A�Ô��z"A2��*̴C�}�&Wd�$�:Ǹ5�dp���n�(�7x?��kȱ��|S�q�9��P�95$�.
��]��0�TB��{��K�C��6��s��2bT[�3GFe�	H7�W@�%�6-AY����lے�Q-=��x���tҲFj�)��
��r��������t%�[)���S�,vߥM��J!�h��[w�=Ծ-�Lή����@#cо� ���PI3��L�>�f��[�eWPu�F媿��C��Ɠ
�3�Ȏ=nt�Tѻ�/����DAh��	���XnH$�EL+V+����m�V=��5��Ѥ�l�����Hܥѭk)��]@�߄9oF�� O��P	�����%�B��u$ ��ML�!�,��� W�K��$�0bX{;i[v'�4A��J�[i�J�ٸ ��LԪ�}W�o�s6�V�n��c��S��3^˖5ב��$���`��Bᬍ�%��(k�*zc�n���[-Ib��l����N�8�S���p���%�JV>8�F�E�]�>�nV�Z%�q4H���J<�8�:~j+���ņ�0�Y�ƯL�?�Ӛ�ҭl�o�:���~c����{��������m�W��9	�fk,�Ē%����槂�"���їˍ����'�p�n8O����en�<N\��/W����Q}���Ji��P��Fn�P�wts�CA�=��3,��MC�2���)>T,��|a��Q��$ڐ�v�ĲF��dKb�����Z~/�M�e��-�bإ!Ġ�Hܭ�l��ɾ�a�8���(W����N�WU�����OL,��n1�YΧ�k�����hϗ���cџ�X>�di���Gy��Z!p�t����z&|a	�m�=3iN�B�cM" ��p'���<��w�KR�1�F����eo���f>���@MhM�G�s�g^��jt��T �&C
�5בT@����E��O�Ucʇ�E9���l�dN�ޥ���kG4����ax'W�v�Ż0P��m͔(9-�p��1���f����Au���dr�c�����\������=�o��w0�˅�h��ps��|�h�@3M	��[+�
��F�4��������-�W��\ �@�G'�q��e;J!���c�s�O���-���"����7m�>����,�t�ֳ�A��X#��j}�}�|��6��v�9�
$�|m,<~�AB8�Z����y�D�C�c���%�U�H����3�"YΝqAAA�x���ƘI�_�ce��4)/�?�s?���l 2�>a��
뮶�G,��e3K�uWqE�&��H�EˎN��A���W���}��L�f�]F�Ŧ	�]F��j��gS��Iyp����j�;<5��5e�X4��V�e����J�{@�V5���W�>9E��YGI�)-��h"OW۳� ����P�M�R㖸���L�I����Dg�2�a��C%�5
�l7��^�q�'Xe��5%�?K���1�/"���}��VB��~���)z�b�f���}9��4�~
*��K�V��d?�*�v���GI��4���	I��I�l}ү~
d�Z�Ǥ�c/��FV�V?�~L�A!��3�Zo��`�fM�	��jp>�=ҩ���=��:ãE#�tmWR��;����/�O�Xz��s��$�Ot_��O�^�5�
��_�w >{Kg;<�� �6�B:VΥ�\�'�9��o=t� ���9x��cޮ�E����mk<�4|5�j�#�s����N��|��u�N�ϰ�, �k����e��\|����sFe�{�A��@�O�,.��Y��Y_3ಙ��D^CN���1o�5�`����Rb�c;�w�ٶ�1���|s�Pﲙ1}M� ş�GΪ�ZtO�E��ȃ��D��O�rl+���	�8H>�r�1�!b)�'J�Q�|S:hMS"�m��Q�"Sj� ۃ��n��ӫ��Y�̺��jf��hS��6R�8��I��Q:�'N�on��^XI�y��خ�g�V{%�Y]��n���<6ץ�ٜn��WQ2};2,���<�n��n��_�h��;�yӟ�k�v�K��蹩�v�l38��e3(�ؠ,LIF���r���ڥ��`���DxQ��ɨ�vݣ�!�l]3ᕘB˰U���!�����\���Z�_B�C:H��[0�[���<j�aF����8��\�1��=�/$"��n�IثY���J���|�N�	fI'��qJ'�A�l�ڗ
.���K9ث��3�CH{�Cc� �G)��K`
���
��n;G�ږ
� W�	�='���`&�diC����~,�Z�'���l�n�I�v���2�n�GLN �����h�^�?N��-4�
�<��bO��2�qZ�ݳ�J�RgJ�%�2�����(���K�'��!��~��a��W��"�*���|���|t�}�0�8s�{��~7~z�#��{晴.��������*���{h;E%}��(�]!�2.�F&����i�J���נ��x�)/N�E����L�����K
����7�,��<�x�K�*����B�X�D Ǎeh�Y���
�FS�"�V)��焅D(z�vÉ�B`�,/�eZ
��ע�Q���r��#g��d��XJ�`�Z�Gc�'.C�5�~�7X������e���{�U��|�:4ن���@
&�]�F����IȞ8�f�Z�Y����M\������j��>��*�25e?�G׀��e�垙���Mf}���W$^��s�AJ3pi��և�p]�(��O�����X	S����]��~��9f`gJ@d��r��t�1#U2P�Dm=�A/e7����@�{�yWI}�LjA�M�e����#_��$�4.؄�m�'%X��E.N{�v��#��AX����u	�2"RN>��#���6�����ss1O\��|�fs�v��"��e�h��`����b�|��B߼��LM�J�wP��-4.
4BF�sߧԗ�$u��$3 ۟i�3��~o���h���t� 3��a��8��Q����߇�܁����Y���N�&΀��A�a`j�Sbn �Ůjs��g���Q��g���j'̟J�n�E��W�t(	�-s��V�0[hl����`4�k:x%E5?u�ϟ�j������<����S"��8�����9�сl�f_�_wT��R�``�f�%9�ZX���ȇ|$�����Ƒ�n-˷�IJ�&SZ狥�]���l�Y8�~HZZ����/md~~E.�������w<�s��|�eK�a:���(뷑q\B�ϪD����	׻Q����E��$�b+/�;E��� �?�x &������ʄ%�Oe�H�EB�����J�Ș�8�Q�,_t��R}6�����I���)8�:�d(�w��cc`2�-���ʳu���#����a���]D�(�KE��T��ٱ�B\�/l}fY2L�v?y����q4�5��OGK�0����Re��s�h�V���5���oz�:�&_��DĲ���4�*R��J�P*#���Mi��;�9�辊�W�9���9��m�H��W=�5k����|^_��C��A���7�n�"|����ʨ�� �Y*�,�!�9fj��,�n�X�p_pj�d7VhA���Ō�� ��K('�D�1�*�+���,��:�d�ʿ��^j�Kf���.��Z�v�9�ce[&<*=I�0h�D�}�ՆM$a�%���,g���%TfD�hh�aW �u�3XJ�n�gB`kR�Q�5~\<̩9����#�'N�ޙ��s�١J/CMܳ����b��f�b;vq�$�W��\0!�Uρ�Z�'���R�%&�<i
P��������rN��ӭ��V�� ,�=m�"� �C��O�������{���.�*����'�4�/�D���Ӥ��P,�H"v�b�K�X�a��d�W^g2 i��ĩCW� |m�D6Cuh�ԝ�^ؖ��ű�ރ�Ps| ���[)�-fƇ��H�<��*��/P�rN������,	�&|���FP ~�^��S��+��>��2b9O����\����JEaB�ˋ���Y�Kr['d�ڜ���(x�?��i�2����?�ez��ĵ���3Z���ʿ���I���'?9Fǈ��i�n����ۮ�<�Ԁ~C�B�Yxw�A6����jMw�*8D��G�Ev��o��x��.��$ce����0�Hʍ〥k6���J)i�|���a��\)*��J1��4b�(*���w�=�EqhM��dW[>&�2��'��jW�Og	Tv�[B�Mh/�(�2u�i&ĺ�
�|�2_3Vg��w�w֒[�9�{��tt��ԠU=�q���`=U�)����̥ڌH����k��%5��ti�WPcSI��L��u���9�� Idh�	��N�WD��%��I�V[����ߴ�z�ҽ���z�E	�j
"�05=M���������E���20!��]+��(q�?�FW+_et-P`��B�Qw c�[�=��8kr\�{�@{?�_@�G�W
�Uw\.�V�F��P���/�ۇ�B����n`��:^N޲��Q.F�͵�đm��ȐK�X���Q��4����HMp���(�m�1���7m���Mr�~���©E�Qt�����-�hW {u��Y�wu���_5C'!��)�L�R�<�;��{�UP��i��\*m���/���r�/>�.�<ʴ��!xGt�
9�"�1z�"���[b�ĮCv:�u�d�f����}�hQ1ݏ|��2��������,X�l{�S�OXC��z�)'~P���_B\����_S��
tl��FJI
@�9i� ��ZGj͋V�B��[h��n.[�ښ��Gn�����ݏZ�d`�J�D�8;�t3�'nǻ�h࠴e�xkV<��0��b��>� ��u�-9��b.�B�Qhz���Or���uܶ.�K�g�8�y�hDr8�L=���-j ��$���,xJi����-a�����;�&��<�O�� o�,}KR;?C���@��a)��o��|�<
�����;�v�+ɹm�}�W���
Vx��V�n���\��-�����T����Ok���h#���j0Q���Ch�w�5���P��fsǩ��� o�*��sQ+WB:�!�� �& w^Jq����r[���_��f#�O/��[�]$�[U��| �L��}E)�K�r߃񂪘<Tf��F!R��������S�.����kI ��>��~j�0;<,Fqt�E
=�������)[Z�����:aco�AH����Y�����[��Kx�d��#e�)쨚��BN�.h;�'R`L���T��?2R~�v���|�w�"��+R�9��r%�{.b9G��԰�5�}������Lr�ԕˁ��O����U�� ��i��9�$�bx�P���V}�e���;-1�~�sa��C�gY�I��Ǐgh�]�<`4�e�B5L�����W�oi-F��~�q�R�B,3�I=�І��'y������A��Yog�.

�l�?�p����ȶ���%X(y��MN�b�1g~\���J#�o�`�;�6V��"eW˄[�&��B��v$� ǂ��cٕ��	�T�_��,ce""&��D�Z?��\��8��~r0 ���HK�k^�nIl܃�9X�I�d�FƜ�f���*
�t'�g\@zQ %��TK�"_�(
]�"�	4�B<�3�U�W��߄�9ΏP�HDa>��v��t� �9YW��O?/h�-�%�Vt�2f�ڕ���N��nH.(r}���4Z�q|.$֞�S	�WD���K �\)�D�����[Tˋ�ᖼ1��W^d|5"
��D��,��5C���Y�u_O� �Lڹ-���_��Ԋj�<�*k�X�V�FMLO0�"���Ʉ[[�92;�נ'_������i$X6pF�s���P��.8���W�s���p/�f���3�e�>¥%�0�<Y=]࿡��'aN�R2��q�
��>��*̠k+!��I�NY�I�%Z�=������Qp�CY�;�2}B����H���yDU��W=��g������Y}Y��������6`gARt*]��^pm��{���z�w�|�THk t�g!`��.[f	����R����x�T���ޒ���~�q�����~#P�V`vb�GN�IP�L�W���g�i�.DՇ9�,�p������n�\t},�<�$d�
��k��s�u��"��m�«��z����K��8q�	}��(jǿvX�	k�m� ��qɌ�b��4��8�m�,Egʀ���3�'�/{�_gZ(�il��_]7B�R��!X
��g�,M�=E{�Ʒ��D���v^1y��P8��I�н&��@�)d��=�x?s�##��fH��6��A6+�	�`eu44�RƆ����ֲ}��P��IX��D�/`$~� h2��Yo�c��?0~J�9���`�Ϛ�v��]�h��[��Nbp�{Ė[L��@�||l�R��:��0��88Vu@ir(��`y�>��J���aq�Ō��&�d}�qqr������{�A�!:�I��o�ǐ���6�n�ԋ�^�k�+����Oi�a��G�-p烿����{ �#a�%xǌ��ay.IS�`,��r����hхD��c��$�(^T���5�~��{hpˑ�Ow;��P�[?#�M�I)������1�z� \{)�p ����S�;bQ%Y�>���ɬ��=���/���̊v�W�&S�X�꿯Oc�=�A�eR�����ǭ�B�޾QΨX#��m	w�:j���Y�h������a:�&mN�C+���w|^��2�J�M�޷���=���?�6xJ��9b/cFzQ�����ْB���pc8B|x�@E1�U�<����
��6�q΢V�(�&�F���6�ݿ;�RR,Z4�W�A��@Ti<�{9�z�g?�T6|�0G���OYo�`zE�����b������uRm)o��ךg��7��\�p}���C��M�AZ<$;�
����1DS_�uUBg�2`2�G�K�����Y�L�Y�
�>����$!S� ��iJ�?{��lr����I��4����7�\�F4Z�f�z��}^X#��g�в2�xm�֖��M����k���sh"B`�G_�
�ӝ6I�b���
r��{s����D���+�O������J~a�pWkjn��o=ɨ�o����j�0��	<>'�!a_� �0va�j g����g�Ƿ�+�	�O���	|o��[�/3�F�L�0 (�b����&$ j��5�k:��}��}5`�	��ٍ��`A�s(O�=ۉb`�T�b{�Y�S�3	�����1��^~���{���c�-������1��
���,x���4���We~�޲	`�k�c2EZI�g~k�.5�
�¸��v�;_9�I��*��,��Cmݞ���h���0h�Zb3n��G�]S��ݷ����g�W4T�����4�fo���+�ߟ��t�( �a�9]!.\�$�k�Q��U:�R'�g�M<�fnקwi"�1�<ز`�$�ŝ0<N�+B�ܫ~�ܻ?���-�.v�`�0R��m|z VN@UI�Z�LqP	乆�	\D�S��p�go�z�
��f*5%�y��;�ɖ���)$�k!��P���s��Z���J�7i���8����H#fu��W�-[�P��ܤ]�n^I���KB����m���ͼÔW뤠���.��e� �oz��c�F�*x�b���7�q���ר��8�u�
X��(�Ү�_C�3� L����u�3����^�N,!�s����'>?�ek?RL�䇪�a-�,���ޑ��?������z�(r/��s
́Vڀ��X�Ffh�bT� �R>��q�4&��%T��P�i7��8�$�"Ӱ' �دz���	�H�-
`OuZ�QI����!tm�9#�2��@
8S��➑ݝD�0i&�y���v�7�V(K����|�k��嚐\p��-�8E:�.{�
J�j���d|�8�^Af��>Ogq��>~|H�黧 ���;o��:M�U���}�S5,84��@Og�@�|��)W4�ڼ�/��Ud-�ݔ-�R��CI�҄�M��mrXsL�qm�X�x6
�s����c��0�]'��-�k�|�K�L�,ɘ�$i}�\�/�ٸ0cEaw�>��tȥ�?=�b6�E�Mɖ9�v�rC1���$0e��oUk�-�p\�#CD����|�}Ej~��&�cl*�^/P$Y����lv��*�d^��6�!�i�w�Ĥpb~�ow��zc��|u�"�6�|�7髀�3�d�����{�/TFG�/�su[ �s��^�N l�hx�'$�C���QTE��PE.l�m~��y��Y�O���nNb^�����̫��m�ˮ̮ȸ,�@�N]��r�*�yJRl+�U5��f��qj�O$��zX�;T
��*=$fG{�@~A���&��۶a+ː3�?�1�4u�,�π&z�XA��#�4���T_��v�H��_-n�=��10&��0�J
x˽���<U�e]�}�XGЧF3u�{
�ތp���H�,�x8��G"��8�97���`�0Q�MKρMf9ypq�I���R��`�4)}�ka�A#�?_n8�.n  i(��<����2�Y�ǎ)e���f�'�ȏ)!6�U����"�8B�s$
$]��Ev��Rr���%b����A��]54iv�u*��1��$��`�x<A�^����/��|�Wn]ݱ`���b��Y����-��Q�2Z���߯�ݔcXx��I���hH/�$���ou'�3�G�r4Ct�K�o�
���E��I��	,�p����$��GeS�;rU�D뚪F���]�Fx�g]��_����a̘up�4i2�D�Q%:����{i�qx�	�/���%�sh���H���*I���9�|L%�=�
��ǜ\1��-��������3�r{�g�Ь���p�������gM�BG�����E}�s�-�K��{T��l���8��v�.�p��X&�ח��$R^�V��<sƼd�Qi�M�Wz�?}v`� �ܽhG�&�o6�V5�"1��n��>���U��<�y��д�P��u�SFt%S��̔�aYz��_E����������Z� -���H��@ۘ�U��G���aU�� ݘ/q2`�o��b��M�۴��$�//yX�A.�'*W˾<I����}��$�_����ڄ�uR���Aص�Q˿(aY���aC=��oD[���TVp��\/��/;Ude;rO�iJ�\2%��� ���X0�ԧ�ArQ�j�1�K��@#ĩ�^E�Ky��}����8qw�o��!A$v���������1��ͩ��9. 1����^���nug.s����eR�l	�h�R���[��K��h%� ���u-�oR�Iܪ�M�i��`lN�p><ΖիAp�@�{ȮO�T�_��as�2��2B�����u}�*��l�;A)/��f���v@��X~Ru��t�0�aB�xA.z�S�>U�Y�gy�w�\iG��0��%-��e�C�ٷ�L�ŘS��~�S<u��$��SK�8�7惼�@�)���y��Z;�և�!�XL�=���x���W���źg|HG�Xf�B]'+���I8�����1��n&���iLr��[u�'�݂����$�D��A�%�)Y���~Wݚ4���� ޑ�A�:G��8q_��<�_0�qXV��FV�����/��ik��<sO�/E�_:/M윫���h��v�@��,JN=b~$�����kte��W����c9t'%���x+�,�u��0y��)!��j���N�c�=9,�`��
{��Aw({����M�����뼷N0���;2�!haDDy������O�;~����Hh#���
��W��V��u�3��!mt�cW�����O
�/������E��ʜ�J+��?�	SX�[��c"�a8���lڴgB��L5���+j�I����AZl`��:(�[��n�o1�G��0���J��:v`�����u�ܾA���.��A���ݿd����p�O�!��s�qO��k@�ed����LM�%�/ހ�֮g�׍DH�x�k�"�A�Ҁe��P:�nsG�Ħk�P��oI��7$��w�&Um�v]���J��k[��f3�%Q�{��/ˍ%�2����y��������|u�4C S ��f5�^�`K���p���t,=��_�GP7������#;��T�KI��)�R���[��8|O���[���,3gO�='NF$��LE�~t�l�����<Ը�X]R�����X/F�K�#vn.��ބ��'CI��Ԍ�tv�0�&&U?�&�u��( �͵k+o�~��4�rHRpwO�cv�#�����0B�/��pD�E#{���<�e0%/���|~(�#x^�h�o��r�u�R��}#��]�K����6��/�(��'w��F3֤�'2ލ�3T��=��;�HhF�i5�.-�/ꌄ4��i38EG��kR����Z|8_��p�D�1��C�<v��0�(/���R�܎T�M�wЬ�MQ�R�l�R��iY�U&����Z|D������-�>j5�.�|o����P�bч��r�x\��o[��cF�*Biie���7V��R��xo��U�]~��P�=C�?�KCpQx[�;ﯻ5Q�og6Mc�l� U����F(f���c���*�g�5�hS�Bp闛�cșC ��5�Ge�͝��y~{K�[X1����@o �c��7�e���q���e"Oj?�݀���${4ɦ�K{�!A�.����Ue��5k%�LV��AbeF�?���Fo��Nn������v����0&Qn{�����G u����s���*R��	|sA�Y����'��=�z.ID���&[��R�<*�)�h��t�?�K�4�Վ�G�}/��2����˃��j�+A�],��&����}6���i��gq�p�3?8���f�f�n�d���Z��܆OF>�� ���A���xkjla�$R������nX]�?�� 'q��L#W5I�tH^�{��AZ1¿L���l۬��T|w���WY���}��[�oϰ s�r�c淝��a���bY�u�9�<S���5��ς�b��)�V fm�UD�xL����{����n�c�n5�^lV_H��Kǵr�0�jE���Ϯ��z_�V���p�9�$-�d*W��@3p��	�\���Y���Y��]���(�G��ln���F#Wk�Y�a+xAOe��0"�?��>�Or 8X��k�eu�y��6�`gK_���Fʤh��z��S�9c.l�4�n�a|���qu|�8��'�6�lM�$X6�0��c�`���_gv-B����R%.	�Yu�e�^r������7�ʝ�?&��#u�
M&F���)Ќ���ZFg���Ai�αl����Df���&���ٵ��->3�b�wZ#A�"��/ˤ�9F��6V���_B��s��}a6�/����	.�}�JHD���r��$Ӊ NL�����j3�YSQ�G�B�첻x	ȇ/�hg2U���w��Zv�R�e�<`m�Ǔr�]�}.W�s��I�%���φ�u�GO7̨���m�ײ��Z��Ĩ����&�`�Ί�����o����7�ڴ�h�z����)����n�����-��U�[O0 (�;�W���MWb�8�K�+�������9��p���Ȕ�`��'YF��9� �i�6�ے���%���.�J�:����0\=�u�.o*�QC:�X�E�`S)>imqCŬ{��E��=�ah�DKS�1h�@�I�	HW��"�;]�w[E�3��~���0��}�c���;y�"bCl4o<�H�:1V~ί����D6��[{��V�0��
6P�כ��Ƃf���-���rd��H��?�9s_�� 3g V���[������1C���چ���<�÷ǹ[2���נ��E��l}�ٛ"�T��Sq�6tM�A�Ai[[�5��~�G�.�� N���eƶ;৖;#��X ,�Ȼ�``���m�h)���t�&� b#�H��s?����E�D��N,�7o�&���yHzNk�� ��yZ�9@�02�;m���I�$�2�^.��>��ܯ���2a�y[0�l7��Q���D
�e+x:�����Ʒ�WHfBq[�,�X�f,���$w��4*w�o�G�)5 ������I��ݨ��(��gmً�I,v�[,��g�T�����Wj�����{l� �['c��=Z4� �W6��ix�����?w�r?}��]nr�ñ��fg߸N�������┠ �����k��~��)1�iK��[�]يw�pп}��x7p`�Z��6�"dw��%a���Y�N�^LLH5�PD�kK�%F��!o�T�m|��prųEf�@+�LM�|�^X��_��x���*����ů!Up�.� Rq�b*�㇍eF7��D�3�i��6����*V��#������`.�h{^
��S���S�-��w�9�ӄ�#f�R�Ҭ���#sgb�?����&��:��:�XF��bxJ�1(���f/롇X;Ω%����}������a1�?>(�c�Ay�q�+Nёx�2z�醥���է'��R��_n�tgC��$��T�KL�e?���Ȫ�+��F�)7�]�X.���m-�ķ�Lr�4H�t�z��,�gFp׿����O����B�[���V��E�Rٶ�(���FY��
����)��@=����G�[J:�ǯ;.V�_��	�0m��A��
?6�^���s���%�������j��~�
@����:�?����H�:��u1�m�z����~:�z�	wY5�(��.;&B��`߳_��271���d���!zR��<��F9��n� �hXg����*p,k���4@Ť�lg��Z���
b�e~I�F�w*a�Q�Y����Ox��7^��j��*��F\��N�W�1����e�}�/��Gw�������WL4d�cR����a1��l
uIV�l��u�گ�W�w�t<�����.z�8�n!��0�� ��ٷ|}���8��`M�@���`j��Osx5�}�{��� ���2m�w�4�+�I����'��Ӵt�U����T+��N��ʴh9�l�D\�5�a��onR�87͙y��Q3��
�*��un�/]W>Gj>9y�X@In�%!�dj.�j�R?�u�v�t�3A� ��6  xU�?��"���"�%��C?ԬHow��N95r�şy�1�<���Bѫ+��;x6�"���S,%-:�A'�]��ey��tG��b�:��F��L7�ѣ{��C*�A/G��;�Y�����mU��Fj*4ҡ+�ͬ��n%F5�"{�)$�Z��M����F̦V��V�߹c�"T����dU-�'~-1e����	@U��R�FL'�.�½x�n�Ua��	�������[|}��.�S����'�S>`0��'�oj?�eU��{$.�KܠU�VT��ܺmUp���G^5�
�gf������9��%<�14I�w���{��L��iƄc��Q�J���L�XJ��cB�<�*,	�㼪�����k{bl���� F�O����U��M�����9O�5bN��Z��&
b�f�ЧˍP�2��
�/b����+�T|p�,�����7��tg���x�뀠kfq'�Kxl�J/�w���)�q)?(zjR^��8��5M��ؕ�x:!;����mO�]m+%��;�4��Z���No�٤�����ϓ��'�S�����H2 ����o���YIM%[}����ٴ��-��D���A*��ړ�q� 9x�Q�/hPB�Ι(���Ixw,���\���.��Yt�>�v��5��=Q�f8|B��< [7H'�=M~B�|��XZ�B\N7�U<u���q���v�ܔ+eywd����~��: rX��:&^�z�LmK30����7a�Z���I��g�[���8əW�(�4!��`XW|��t(� f����&{:k㷙�iɣ�6��{dS^�i�n*ڎ�+����L�Y���X���>,9&�/�n�M�����
�Ջ���q�0�GZ1��#�/�܀t#{�՛����=S�YwB΂5�[��/Z@����KFwn(�۪�ކ�A�!��|s��k�aԷ�0���M1��"�_^=<C�b_^�i
͈��^�=��l��C��1E����!-Z���r���.��&�g��/��)�����3�Ll���w�q|X�Ӏkrነ��X/�.�LD ����W`��-m��eH%��������d́�'�����urHs31�C�E����
/�a6���
MP��h�R� c7$�5ʲJ#f	Nh�c������gYǏ�!����;�h�`�M��>�ocoދ��2F���r�d#��>ف��	��R�2ֿ��S,7�ܪF�&�RQ^���4.w~KA��b;�*_86�Xr�G��<��݃с&�90�G�a��Hfi�el�qjW49�39�
�uD�$Ty�����L�eb�2�qB6�0�6�ļ]�mZ����nj"W�m�y���u4� ��ST������c�M�dΞ·,�c�
{V��_���?+�����$���j$��N����	P5L �]v��*m���m��}-9.��d|���-3�:���P~_��{��������5|�� y<����!0F㣑Y\\��p�Ҝ2���_,iƞPr=���j �h��]�� ��h/����8;Y���f�����j�wbf������(�a��P����G>�B�ws�c�	Sj:�zd����	�鬻��)�_ۯ�\脴}�>=�Q�5����K�����NŷtH��ɚ�C$.PE���DU���&��Բjt1O��"�F9G�KR�6�&����Zu���RRg�O�����P��w�8������^d���P�͏sH��H�-�A�c��{�+�i6�޼o^Tj�OWI�Ȝ���դ���4��bT��T��Ĭ*u�a֤�瀊 �Jh�fK�l4D��6����6	蟺F^u챫�D񲅾x�U��<EĢ�5�y"*�B{?*8�i�{�>X�+d��,��ю�gJ$�%P�i3�NRŶ��PQ���3J?0��C���{)Ø�28�f�Q5�u��t��^�*װ��[�@!�z�/�*�<��5x�P���x6f;�Q��Oi�Y�@4|��HC��kT��'�tma9����]�e�~E���r*�&M�β���]D*R���h�����|��_Y����>�H3�pU�d��`*�'dW����`��,���ۑ�(��U�-�����}�ܴ|��e�{�|緳Uq��[�L}����<�%���h��zC�	˶�I@��j�~�&R%s�6�y�t[,,�Kx�f��zB������q�&Q�M̬c���L՚A��m��}����*{��x�h����I���sr1�̥>}m���H9����
D�%�k�X�9ߦy���V�e����N�<�X*�,��%m��`ķέ�7܆�����x-27[�%a�_o�� ]��~��K��SJf:`z�"	Q �S_�f��O��O)�A$��o��s���E�ȫn�<[�F��U{h���>|�s,*瑟�I��kФ����̼z�R�,ΎI�,�A�N��f2"�<�
Аzj���ƫ��^�����+��W�0O��� ,
�)��܁��=�K�!����t��c�	��g)"�޽T����k���L|�9�o�T;�u�KنV��ueQt R'��ʹ��nPe(����]��M7�,��u/���|%�eR���L��<����H<���G�����q�c46@�x��c$��fv���r������QO�EO���+�Z��囪��q߻0�բ�db�#+�|�eiJ���3�����t���B1�֑b�Ig���@ï�7�h܊��Θ���@$�w��z�o֟�u��`�o-�L�B�g�g�
�@I+�����g�~M�I�N� @\��ӫ!o]�~�&���)�\]GeL=;�>���.ƹC@jMI��q�jb�����r�ɱ't��ݘyyu� \j`����_,�G�6$��M�ǲ�;w������q3'G�|�(޺X�"����dB-��C/(��9�7�L��f�úK!����6�_��<���Xc�Щ+0��~���UI�!�s�a-Z���F���=����/�s�Q�$9��� �\�$t#��L}��|3/�1��`q���6	a-%K�"-�����e���#���@��Pz����i���-�I]e��O�R�}�pB��G~PEad�d�-��[�)r���.	�6��,��9o($GXϞ>(�*D�=�������?3դ{Xe�m%r#�M�]�n*�[�|����}L^��b]B �P@��C8V�$�!�8���rwmR+������lǲ��|���iO�2Rj@�8���+�7h����ʭ{�F��V!!o>�oE��	݇��Q;��	��>��+�z��'�:S�ɯ�ђ9Va����V��^.�u�R�8�}h:�\��2����轣�m���	�sK�2P��#�P^��Bg�Mʄ�a�Z�uv�2�Y�.6���=�|���M���ˍ��'dF�>�ľlPԨ��5��S�GԱ�K�, <�r11m���G�&
&>�����yPJ���`9ORڛܐ�A\n[z�J����#�+%/j���Z�5/a�k�_O;D������Q��s�\/\��͂	�곡�eqHj��t�J��^j��Y�����0��p�ha$�d�/�fN&W�ei�-�3p��x}��7��ߘ�M�����	u\�O�;z�)@i��芐k39g	WB�|E ��;B�P1�>�|z�^�75a��U�iO
l�)t�̺=L�i�j։�]��M+�HSbQK�9�O 
�#�>�
k@XcwR�A��]|�ƫ�3��/cK��5�/z;��mʡ����m�K~2��y��?G(f���J.s�q�k�%� ��r�}�e�K"�57U� �tW�m	��/�������#/����g쐊�TQ������&P�y�M��H@�3�="����l	���Fem�K���˃B��Kc�#�*�ɇo[�[ţ����P��Aq�So���T��7��#��7yn����]pؿ�e�hQ���z\Fޚ���@����,�ճ���(����ǧ��}Cԕ�?���O+������[���m�������#��H�9�^rB0˖t����+c��*�`��a`������!��`�O��q��/���и�+��Q̡U�[�����|ѓD��2	���H7h�ˡ9�NCы��ja����^:�-�N��M��F3�]��߯�3L;*X�k;\@I��>��b^�bV4�hlr���6 =�^4�F�-���#��Z���Eg�,��!������JO�O	��=A`�Hx��3�l�>��}�b��%mUE�#s05�7,�����=&u�b������ʌgn0J81e��Yo�P^��QQ�_���HveM���X_1�,tn�ޞ�M|v�? �]r����~���d�S�.�]���۸��ϓ���K�yBaH+���h�û�%ղ@�6��w�q��}�.)ƨOw��19��Hf��nAtܖ�`�_�z�9�'������{̓l3��/aЈ�vg���d�=:zT e��@����-��,�.�d�iY�أ,��[7c-]�zX���Zb]���)笛A�ߕZ//��rJ�͍oTol�ۨ气'�2�͂cU��#ጶOG~��dPP������Q�R�Xy��ʫO̜�X^��r����^��Cv��[��'\�;&�ghf��t*��I��Ɩb ��Jǭ�x�o l�z��ދ��E��r�WJ�mؒ�v.� ;:,�)�X2��=U	&NH˥������W���< ��ւmbY� �y�jW����߇N�s����?Җ��x��|�z�-��@��0{�fu|��x<�붭#�	e�DeW�&|�<ET6�[���p���`��6I��Y�·��؂c�&��l1����]�G�p��Z������VҖ�g��яL��`��i5�
ӯS9�5��M��m=>=�Ɓ�5LB���m]�(c��մ����N�'�=�Qۀ'�����Ԇx+����>$����7{6�í��`��.o�/X��v�qM}���w��Or���������79z{�e�!��i��/'(�$��E[j�g�P��0�T��C����[H�hq1s��U��̪q�.���p��s��65�U�d>=pjo}�
��+o�u�.�Y̜��7���w�дf���w*��P %�$e���P���(c/�i$ĳ���>�|������^uc�UYN5�Jj���v�[���JmfBcg-�,��&�!�TY�!ej�����0��ԃ��U�~�����C��S�D_�
�;Z Z�@O�h ͣ��9	Sևǔm�{+
$m�����˿\�������T x{����-��V��Q�����:#�BMƏc����V���fu�Iʎ=UGUT���uue�.yςF~R*���T+���Tjz�Ci7l��Y�����E���֝;��vVU��и'V�& M��*,+�FJk)uK@a����'�շ=���e���&�"ґ#�~z����6��'+��=
a�� K$q�u<�7UhT�p�oLΟWj!���/��r��ɒB�����+�9�M��5>�=����8\����2�T�>�D�!ʲ�;e��<)6�s�*�5�m�����z���Ww[�#�[�8ӄ'�X�	�Dr�B* �!�J���40��
�]��eN%5ǩ�
�'�2}� �9���%��M��������#G�msU5�o�\���N�#�?�{![��7���l���d���s��F�TW�٦���� WX�~ӄ>{�H�R��ѡ�>��/�  ��ų��]P� 	L�Ǹ[�Λ=xL^�d�4�K7�OQ�p ��"i5��A�����m���2�����;�"^����mt���@���Y�jN �ׯ���a�+�`$L��|��nlD�1�� g��.!���%���I�A|fY��ë���͖J����b>dW�L��ࢹ��\��Q�
�*f!!2aُ���`��#J�qJ�*�hDމ��mS^��_��j}��-뉋6D�
mvj�I�DZ��9�nt�U�}ߟҎ�?v�	0��~U�9S�
��[Q��P������"҃���c�da 3��������������ښ�=�o�u���MVC_�(篽�8�Y�p�;,�Q����t���U�3��s�����=�80�"�G�M6�S�iX\����G���<Q�e\���і4Ύ>�*�z}�L��V�x�7:c�����g�QC�O�oM���$�L�����8�61��{��s5�V�C�=�������{�k��;��U��!��v:����)��0@yS
"�D��Ϭ�����;=�����t��M{��TH����rn�&qk����9��Z̍����Xp*x��S���N!�_�06�R�|(&5b)�4����[;�.0�m��i��Ri�׊������4Q��<�R��,���/QK�b�1/Tz8SO6�q�3Wr��;�Y<\X4Ԭ���]���)���q1�'2��x%�qv�4m["�Z��?���'C.m��ْ��,��썓[��5K�jR��Ɔ�����7�G�	c��?�,�+���n��x@��IK�v�`L_�(�hy��Ƚ�S=�߯��5AX�&����j����BV���M���P��_o��Π�Po]�7:����^'�p�O*:�h�5E�B�v�0<����*�{Ǹ��?�%��%�GJ�JÞT����{�$�U"����B�5�Q� �/�A�@��e��1��!(�)���Ҳ�|2���u�oǥ�$ҼO�*1��w����~�����H��v6?<��NJT&ݪ���W#��#��=b���t�ۂGO���Uq��4��V׸<?ԐXfaYq��v�ۣ��ԗ�+\���9lC灶�Fo�cA~L�7� ���)`����+ ::��t�g�}se�/�^�a�s?9R���֏/�=�C�Fʵ�Y`�W?=#�%��:�������?�R$m�jG�3�����pI���
=��(YUm�v�M�C}B5Ƿ��4_�PT֬��i�C��iP�$����a7R��>p��hۆ����F:]o�@=��5`��V�ϴ�Uv�� ��"�:d���QS�+p
.�$��*�� �`�z�����K������)�8� ��0\i�����'��-Ɇ�K�ShܗU��A�"��W�^��VH��Q3��/�8���-�u/O���e�*5���T*ņ��_���p҉����L�P���
��W.�����;��ǔ;' �3(�//�;J�9$�����T|e�!|�%Ó�h�(>�Q����Az;)X�U��z������*������YK���4^���ͷvp�ޜ��"�To���̽�9�-X0�-p?&d�T]�B���@+��QÌ�M���J�}0l�?,Ȧ�c�
�2�jE�W�����L�.�����
�T�o/w��.f]��qA���
�����U�[��v㍔�"�Eb<#�v�])��Yg'A<)gU���ܴ̯ PH�$
JgT3[��F-��+IJv�����`�A���3فy��߁��U�� �*Эg�XO��V㪉�&��XQE�t��?�G�o��Ai�$�����]H��ΚK���:��@�~�);9}�m�o�OJL���VK�NcFƨ����K��X0f}�2r��$/" ��\�b�#�NȰX~�~p�Xa�	� ��8�2�OЙ����2]�� �4We�E��ׁ�D2
�в D�4y/��e� �{	�N��s�OqϛV/ζˍ���sE�D|�i���"_�F�Ul֊Kc�Y@���3ҝ�E�+�y�/>���n�F���$^O3�B'5Z��Xe�l��MkCF�m�lz��y��d����C�k��S�S���XC)?����"ԥ�j�B�;!�<��f樳6�H��.�k��^7#�I�ɴ��b[���[_��&���������ʶݱ9hmA�nl��������H�*��4��@��7��z~��+��䗙����T��Tm��dW��`�PR��ۨ f�b�qI���I��m]�B�Q��G�R^p�#�2�c�ɓ�_��X  �2��L�<��'�����h-q�Y�#��mJ�9�h�=W�D��ybmL�9��.-�Рf A���Ö:�#nh�G=���Ni�	.�����h�>Ȑ�����IF�N�)ё�9V�+��3����)�%�f�a8�Df�O����� 94��6̶���F!~� g �d����!؂w8.����q�P�f��4�����4X�MI��#F�c���^'|A	f�y�.���֙��Ȓi�)-5�KU��>��V$��E�d�y��+��:K��h\�魜a�m��}}.�j�B�~Fn��~f��;7N���6��:	<Q�+|�A�Z�F��|&�<Ie�2���-���u�������۝�B�uJ���̇&o�aߠ��}�1/�Ku/�x
g/�n�<�(�2��� ���!��~Z�Z��A�i$��<�ö\�cԎQ����?=�l�pD@?=�D8���ʙ���x�?���i�J�VR(_���\.2�����e9@u!7e���ۥ)ed#��z�V
��& +�K���b���]��c�~M鼅��@n���fq+��g�Z�	�!t���MK�t�:�����GAc{�@����0�`��~���[zT���|�2�����A��ф�'6��W�1�&G��#_3�s6ĵ�$�%�V��� ���w�x����n�sş�ݹ��5]Ҩ����+����؉R��K���Q�#r�ck����,�O���)�Nٗy���fFy��
@ 9p�C$�-���%j�|�����=�<�U�+�����8��
�'�,��&O���!4�#�F�B���_�f
A��g������vls~���sK���ڽ��D���ǒR
y��G����F�����[�>z$ea��3�9Q��n �Ɩ�+@��\�a�a��f[��N�-5�0���)��/�%�Epб���N�1:��P[��Y$��*G�DIpvpQ�+'�ӬTo�+@�s\�?2�R z��~�8�=�NP,�+��"����'iU*cA� Q�/3*�za�4��^����]S��H4��H���_ݸ�.���`�}R��R��X���դ���z�d
��M��3_S�������0�Y6���^N˚����x��N`[��+��<�-��k���x�6"��r�K�n7��(8
T�G*{��v���y�����!��X�)��+�V|������5��t���\���u�,��M�=5���_0h��>օf)��Xʋ��j��w����� �u���=�	��J A#M��MԩF4h�>�Ft��hl�nf�ٽ����ˉ61�*L�t�IG�/�[�R�x��(�u~��m���� �Y$�
Ԛ�Ku<��<�F���]ؐj
�������E[�T�/i�2XO��,yrhe���b����e����q����0,�xA:��|"E���b���`W��v��2a_���|�*qHJ&8*/$�C�r���!?��t�T��⑙���l�C�E'6�~�m�2�j��T��8Fa׻&�cy>&K�|Й�hsl�Bp�g�<���(�'�EP/�H��d;��6OӇ�,؄��+�4��䳎��V��ې͕��L���dG�4��S؝n^���؜�T���qD��|6^��r��� �mE��?k�k������CRZ�f�݉$j4���d^�s;0=�� ��ʑ|�WA5 !���(�ƠZ��! ][He��eu|Z9��V|��e�����a簇��cF���%����h�&!Z�V���N���w�O��Vx{�	�6Րk�����rb�q�;�2ܰ��K$o)i�$��y[[�
~X�Cp��>�d\]Œ��}2?�L%	c��3^����`��ZC)�4��iK$����2"ٱ�;k�fWƧ�=T��D/��G����x�LΛp����,�L�q�/�Lř��[|B�@1��u�� �4�?����M9���+����f�.)i�g�㶅���
	ٰ� �{h>_��y));�jY�&�P�e�AB3X�3��9��V'"��a�-�bzz|I	yV�d�j�br��`����GJ|	���9�aCK6=x�m؇�DBm�Q���Z�G��)�������d�av���yG�8��;"�T7ե(��-�,��ǽ~�F	�\�M�aD{s�b��-�����a�<�S������U��X����V0��7S����"bt�E#L�m%+Bl�4�N�I��Y|vp�?X�!�g4f?�(���tR��w^��Q�>����l��T�u$H��wɑ��
��x>@y.u8L�E��8ɴ�<�xuc.w e�%I�	�����k%���T���tc�B���"K%�T[u����:�������TZ/��RWK�+�@�K�s���j�xe�zvn	��q�k��U~c��p�S5�e@=EX�j��O�iD7�Y��ɯ��)��C�'�-F��s���ZThVǼ펇�ZZ��0/]C&��cTHD�����H�'�1����o~z=*�X�n�������:�1�7��/U��/F��p���)!����/B�t��Eз%k31����eh�n�a��u�\�L���2-�5�C<�w��e������?�5Y�I�ֹ��Va�zǩ�B��:jp�m���Q�sл�_�FBP���rbV��:�,�!��K�(�RF�����l��]O��tʓ�3�� �"�5Pjt(�wB��~��Ek���u���
�E����Lw�LۋS˹��Z=@Q�m)�6X$�������D��$��j>�;o�-8ӭF�cy�x�0
��nUn9^��O�=]�s�Gf�G
�28j����0���Q�(±����F<ߖz��H�����0����`���j8k�Kj���=H��߇��R�U���*��Rx?B�GԺ��=)w�uvb8j�.��rBf�bᠻ|Č2Df.���)�d������� �#�����7}Qb �gO_��-� k��rβG;"Z��O�6����^�l
 $�XA���GW�}T/�!�	d��:G3/�� ��c̬ C�ֶ�bc�'-M��x��	�U����li�t�Fʢ��w�L��EQ@	����?�r�'w�2���hU�w,�x�(ƀ������C@7Ng^�Ӕ��WS	R\~wę!��BM��$f�'�*�S�n��{Ll#mf�r�	y�i\��N+�f�6D �=:e�R~I��vd��U�5{��9�iQ�R��*��-�C�.�h��ÿ��E�ܯYb�&��<X�!6���S��
fjOG��߂���[�km�T�(�,sK�V�;���Z��Q!G�0J�, ���Ȍ7�*M��N�&��`'�c�@c����h�=��� ���� ��:j�ɮ<�����9 �j�+�)�ι��
����.�_'^�%��ę�m1���1?����D8$X?l��ا��H��,5�%��9��m��),��}QS�����ɈR��x�#_N܎�]lږA�u�OD�)c�-�7`$D���d�}���#�ޓW�h<��d?բ�j��:�y�P�a�q�gt��\����dgȂl98RzJ����"@���ΑО}il�	�SX�A�
w��`0��W�6�[��1����'��ٲ������V��s3�+�C�W��8�1��������}:j��"�M����9�o����]:�|�ثJm�`ѐ8�sXW5�9'�@�N�	���l��Y���C�گ]��܆��Z�a� ��+n&6�6 ���N��ط��B+�#�B��=V���
�����Ő*ƌ�7ʁ�U��7p{�����2ej�~]P��T���a����ꅜų�DEr�L�":����V:��.�;KR�Y�L�^�	���nɮ�Y�� �fl���`>}"��tc ��mɽp����U����8`�l�އ��g���	DE�|�]Y���5��5�8/"f\���kw��cr�9v&�Tb�ˬ$��,�po�{TW!��b�B�V���-��	�a�q7��%���ť�DP2z�wJ�!.��ܠF�?Q������� �\��b�X��!Z� dS�8�������ۥ���
�3-ｏW�k�z��n��)�v��vw3Z�g'2_cB��;������N�w ��LH�%c��XJ&e�lL�FN�WГ ����<[$i�Ce��g7��xp��U����q�Y�����[2Թ��t+w���w�ӈ��M��N�-��싗f�}σ����[��A#��L��9��+�2��L�yp���Ug7L>b�Dc�����|�hYM�Fސ�ϟ���>B!r������la!�|X+�sB�13
��f��7��(�T��@B3.p|O�`ةT2���M����`��}��x��JdS�W�Q��)�j��r8$8�O�m��W��"�h�8�\�L�"]&r�(�d��YJۀ%o��-$��rJge��b�l<�L� h���yWY��#�|Q`��9�-��bo��A�!��G�n~*�\�Q�/��d ��^RF�?���I�����>�h�3%%n4Ȍw'rđ��SVr��VY��H}����{�}W�PDXW3MS����l���1�]+��m���c^��j�^��1�U?X.E#/�$��$kq����OH)�{mhN��tN�ۖ�&���O�xZ"9x��[d�����yB��x꫗�q����@�d��oP�1�I�v}��D�7L����6`;0I��1�Õ'7��gx'�[�N��p�B;h��L�N�9s.��T�C}�(�Q� z�^�ِ�F[s��B7s7�cN��aE�@���A0h*�2���j��Dw)���Ye�,yٗvؓ �r�a�0�Vd��e��+9��X��I�<����S��qZ��/��k�W����8�b�;Y��5�5!EJ�~��C��7_v�[ݦ��צ�7�~��@���AS'��Y��'��[|!���ھ����8$�^�n���Ξ��V3}��bu��~ky���f�@l7ԑz����]��d�)�?�Ł��%\;��i؅6o�MU���yf�$!�8��A�|U��I<�!j��@�|^��f�9�!��;����`�g�_� �=�)���+}����B��AKT�)���T�	ցTɥSJQ���u��!�c8F�%$��H��E]�P0�3K�+�6�?�x��%g��*�#�7��%$��>�flװ�-*Se�hC����KՍ�t��n�ZS~�H��[Em�a5lAEƽ��g�§�9���n�~�rY����< �>�����d�/ꉪ��g��<{/���g~X�j/^ �!*n%���J��l���p�dH/+p.�'P��f���"S"�W���ua>:nP&�4䵶�T�	Aǀv�-�3lC2�)%|x2�IE��D�XX��	����ڸu�w��X^f��g���c�_o��;Dm�Ҡ��=ͯ��`�3��AdhN�z mw��m�M�f�����`�ߒ�$��-�"l����Y�N0	mO��e U����^��B�ɚ9���^��d�5�&�=�)��R��ǍxF}��M#霻����C�8ry�3��^���Ii��]iV"K �-& $��Qå�U�H6�����k�����Xd=J<���l�����n�V�lXM�k����u�����IBT�����lʉ��Gh��c�[��h��H|]�J�=�EyD���Ͱ�bC����B-fbQD���"�ms��cYHQ���w�H9��`Y͗��4ĳ�+��P��p72
�kQ	W��r
 j���3�ב+_��I��fV/�N7�#Ԫy�9DŻ���2MS���b�{�j���A8���M��ؔ%s�ઁD�y�`i��s�ܠ6,n���T��Vhn�Q��U����O@܍3���/��@�P\�#.QX�(�M)9y���#�x�Eih�di`�����%���T�W�h;L�����:a�!�G��ͣX|{8��<{+^X,����{�JV&`Ѓ&Mȑ"~[Z����Ex�_	 I�od}\�c��Ҟ4K�Akl~����q�9gbx]��D�HD�*�c�����8M�d��Txw�7]�6�ġS����0�4ޝ|�ó��?P�=���:^�{��̮LI]�y�A����^���a?]��.Y���U��фt��UK���u�Q)��4
�S'1�`s[��)�=�s�܀�'Y;��K��U�l��d��j�dM�b�"K���}�/v���niQ�%��8�d�o�0J�|�N0���;p�J���G4q�	(� ��Τ��4�T����=/�J��}M(���� <���&}���a�,�Q^|�D��)Y@2��V����������o*�u�7�r���K�:�߅5�]�����W>ܦ��0�ܺ���M8� ���	�^b��Å@9�􍯷�h�c�L�)-�$==��_J�>{[.��p�:W't6,��!���
`����ʠ���9������gz��kFC�Q_<.���)�#���a�AG��(Cğ$��f)�����
i�pQ�����/��IQ��eM��T��7O��C08u�~��HR=��Z(�z����)O%�����j�_����pp]�Ue��`-�'���K��Ng��;�̽[e��<I�g2z�=�l��K�T�̂�!��1��`sG�|.[؁o�O�P�����N�@�`���~��u-�u�.ټ?z���8������C��5����AT)�k�`ޱ�b����꜖־��*e{���^�QZ
�h90�b�ģ�Z�̔��[wB�e�J(�מ.OH��,4�!��y�A0-e�rH4�h�Q��&�9x�����$���>�u��,�r�lr�`2����s�,[�8�J�])Į�눩�	����HI�9����)��0�v��}�aD� �SxY�Ϋإt;�Vh�"B
�c{�Ӫ�6]U�^���.��]���h��V$i�7W�qt �d����8��eYg�m4*U����:��'�ۊ�xM�#��jI�7;�K{P���*%�\��W'%o��P�;(���&F>(�
�<�w>se6��C�CL�x2��J&v���|n�8g�q��t��Ox��т�}o���#L��P��1$f���̔W�����fH���@E9G,��[���zŷ�b�c����h�p���06\{�{���:�ɷ!��
r5�B�MB��;��<�E��\������/��t�R��gN�����v4#���>�؝�W��'���AL�I��7�^�m%b����CP���7:��)k� NL�����N�qm�晹`��BS6���,�Fa��_r�Z^I�A'Ȯ�R�ɧ� ��Wt��P"?O�d�h�H��D�V�3�Y���v��~x��S5���cR�1i���j��3�`jmӁ>��	�g��|H�� ǂE�8��1�fO\w:�"<h��ˌ1�{�	�6p�w7�Ύb�(g�f+4���ޮ�츓�G�����i�`��1�Ȧx|ړi��Kw��迉/w�i����)4��D!8�D+sK�����X]�)Lűa�����n�u��(�#��(�XD����!�S�!ײ�5��9�Cͬ��{�Hq;��?`���`����8�{�J<��`�<���{���;���!�۩���6^`)���.Ϊ��+ЋY��p��o����_)�gE��0I�dûp	���b� ߺ#߅ߊ���"к"��2#�}M�Q��]��:��)b&<�o�u�~��
��p�i��\S�_??Pq%�=�8������5Uh�5�}��,U���?Yb�ݲ�)d��rҔ�Y]6�� �������8��{�lV�:�M�N��%ߖ~���`�uh�N�yز�C�L �j�JM3�v� �b�f�oi}-���>�Cg��?b~�\���WtG�99��#�Q(���$4��5`�Z����+�H|vU<i|Q��E���Ĥ�ℯ�]U�g͈� J"����Uɴ�J�-��2}�?�l��,,<��y����1`�E]/`�w��X=��tv�K���&�/���z���62�&�Y>-A�Ų���o-�D��0�p�
��W�EO;=7�`����jjF��vޤ��W�t�4����ӕrq�?�>ip?taI@�W�a��Ehܾp�&���}k��㫿)ݚ�ǯp���7��rk^�Ãh��PbV�(�/�B�=���癩}R�Ĵ��8���]H��k1��_�o�+ߪ��S���B�=�e/씸w�*s���B+,˃V���%����yz�F}=`�r� GZE]�}�X����օ��9��Ȗ�"��#�Sȇhѹ�M�V�Ҁ�	�>�Mx�{rF�틈���p�2���S���˦ڨ��әo�բ��]ɤ!)��5|ygEd�.z�5C�:¦� ��̯T9�F�� -�8����������o��0L��d��TpܧĎB�J���KD�����ue�X�z8���({gs�)��iw+t�voV�Y��i�G�8K�d16C`AH��`f���,�X��%��M��`w�>���{r? Hcvc��`��y�W[�h5�dɴ?%M�^��̓v�pG*A{�	�]��]�(�B��#��,*HK!dj�z��	��Q�P�pZ(�F�7���)�K����`E/���@�I=S-���y����͒z�Vst͒ �0) i8}��K�b	a�χ�ZɎMC��'̌��/����Zk��uOp�Z ��W�D-�h
��tuђlf�e��m���g�o_d-H�rs�I�l2f�zjJ�'�Z���=��
��՞���w���ʠR|#�o��w
�&|�Þ�c�j��.+�f�Dt
��V���Z���f�,�]��ܒ��:�r�^���t[�G
'XTI�I���	y�n����A�V'�On̫k����7�꺩��7�lW���H�c����uW��H)Y����d�/�\̭��G�g�b���Ĭ�!��#����!{u�{��sjU�P��b\���X�G8����>�=.MdN�a���ș�)�=$w�!j^��0�"߀f���=B{.a�o��0����Z:x�S���݊�� 6eJ�BO~QL��d�i2�HY��d�s����T.z8�_��O����q�յ-V��*ʹ������j�\[�2g|���>A+�B��?�1͋?r�I����8�=B��^)6���_>�������`7��'�� P�ˀ��sQ�0�l�Av�0@'А�/EpRc���ݛ����(��E̟��w��i��)�nI�%����n�o�H���p�'~�,��a�5�ڟ����N�_(w�����^	��N}� ����
���p��\�����7�3X�kdYd�c��845�n/Sop�?~(M��փgoе�E�լ����/99�LA.���k���n$�Y�|�H�K-E�T�+���߆�ϰm*�k��Ĳ����FB�����alӊ���	r�jh�ת��Z�&�t�o�!���zb�	��	������m�8SϿq��#����~A��L1���:�}߀����(�G���a� [����Z��$_X$�;�z��ҝO-��y��.�|7$c�$�o�S�R�(�j�E1o;��3+BO�R�����U���=�p���D4�~#\Y����W��'�G� ���9h��Ȗ��wj#sB�Z�s�jeX��k�{�G�X#�X�I���������5����k
S�����q��W-���B�֭�k0�1�9��?�)��p��F�[t��s���'��y	�%�f��k�� �_Kւ���$P}Ȗ~��D����l7�	��w�j��'�$X/u�3MT��U.��t�Y-ia�]�wq[ţ;K����5���W��m�K=�Lc �����W:���q���1��J��<6^���-���6O��o��3#�y��[;��/�	��0b�,�l�� �G}���(��hcg�[#��u�g����|�O:�����/���Ę��%��Q �zZ�"t�Ӝk��HNF��&P!'E�@.a����cA��z��'pi	=�-{��}�Xb��[��i$�I���u�.��5��F�h����ZR�&�ip���J��}�8��W�Wx&-vջ5(ְq����Yel��;��=�A]"H5ϴM��5�:CtR���jw�����7 I@.����e^XJ�O�L��1��Ot,�Md�ɨ�&�H2m��CB`~�I��(��V��*��v_)��
Q[U�n5rp��Tr��t�SYl��$Ql�	W�2�q2x�]F�����[Z���*��[sH��e����,�H�,�G8�h�U�Oq���3�ė�m	�&��p�������^wH0Č������i�K�)]KN8y�a�q?Z���i�`��N�?sI߆P�p��.}C�������L6�l{�V������GҚ�P�尊ti�j���3��P��_#���yw��� A99��*���� ,x|�J;�MgZЬ!]���<�=u�"�я�#7_5wh��4=<&���3�`W� ��V�{�,�E�����|�B����1NO��@mc.�T��(��ӵ��^�������#�<\K[ǱR���}�eW�c��1)��o�4�]�Dմ]��F
e���SMdPdl%T�@�Lz��S��9�����웉�Z���� ��H( ��g�w�b;�G��c>�J�r^�:�}����W�G%�~|�!9�=��fk����,��<��ЙҴ���3�]��z2�zfٲ�p��n�S	�

(�gG��Ep����t�<�ï�;��#y�y�喈��G���%��/��*��ïP�y?�����
A��A���G�'ss�=|�#����<��3��$/)2�@:��;a2~x�X-��u�F���F�	?:��Q���L�4N>E���^q���W�P|>{礻��8x,�ԏ�p�]!��ϟT��F� �Y�O�)�K<���	+b����
��R;���וg���a�Ѳ�@���%������T�.F�6x�'��p�y�6�77S�g-��z��a���};%�1 8X�`��Yͥ���~�7��qM�Ի����K�5�$�%�B�B�x,���A��=DĐ���.���Z̊�Z�$L��c�vvF�qeF��v-���
18���9��!e��v���m���n��(ӇW�%�MF�A����X�0R�O��r���7�E��𛢟���Sv�f>%kU�,���↛a��{�:��Es�b�
�q��&N����.��RK`^`\�:h
.ɹ��6���#q(�+Gǵci:/Ӂ���	m�4n� B� ���5^�$76��r�)?��FA=d��NT�w�e Z�-�QR{�fX�#�9fu��i�B�J�'�����2!����+�zx�M�Gd�C�3�_�s���!߱�Z��D-K�2�P�6B��$<���u�+Ix>�/�vLN��'G�|kE���Ge^!�wB1��%\]���X q�|0��<E$���P��Ǒk�8nMw�賱� WoMHʘ٬h��򦢟�Ml�XE>�	=�ݺ^��G��.��5S�ڽ���<֩��� ]{V*i���%�UP~}�2S|�ə?���Wt����<'��`c/"��p���#�"+����>_B � !D����M��XY±��7;N�̆���fWxpE#J���+�j�. |9E�b��A%���X3���Z�_}V����S�v�u����Y��3wӼ^�?�W��,>����D�E ���
1���� "t��������(s�ȴR9�{�Ue$AJ�0�&f%�"����^Ix仙��6\���k��`+-J8BI�CW;@5�T(����@n{�@f�N��Ϫ<h`��x%���Oy\/� U�����3��(��9 �E��?�cK���*���+6A;�3�9:������_��gS����0�z���S����[�I��y`�=t�E�ɮ��`��'��L�U?���賔� p�����v�U��<F����b,�.���n��5p���<�:�&z���:X�J��������B� (tcb$�U����r������;"�^���a@�7���N��l�[���[`Q_��V�4�M��@��n�sܰ�k�Yd ;�I�7P�t@?y<?��©VXdQ[�d���_��U4a�g(�-i2(N*-`���;�%|cV��~D-��?Fz�QE��G"�k��L,J<��j3.{�-`�R�p����5?:k�k5�[vZRܧ��K�l���E�� �X���<��{˳����L'1�����#�eB��3S�t��/"�*�o���@�n�bw2�7e)�w�av���X>j�[�ΚE �w�-7 ��e�(~ q���6��Q-��tq��}SQFK�W���Q#�8�D�'H,�=E3-��F�����H�.�k��>���ξy�s.����N�C�x�2������]&��VNaYj�M\fE�6�s�bX�+/�ɉ�i)S��g\\K�] ��b0��/z@�v��p�Ya-_���_���%n�Ӛ�&��r؅#0��%V��e�v�o��f��Kfe�Ë�É3�*hm�$�*/^M����� ���̲��>�22�i���I���v���}�D4;g��=�Tx �e��.g�G[��L̋��鱭�N�;n�	R��2;���h�r�/�'I�3�dJ����L��Q�ID^�0r	9s��oÛ? \�-Z����BO������J��t4�̭�ݹ�UIn#��1FR����w9C6Q�ӐKHK�#��B���,�:n!r�qbǞ�6ũ68p~Y�sv���?�Hߓ�Lht��m_�?_^Ο����(J5��G,�W|KU�b�ra
v0�\9\�A#$�9a���[�Iq�<��V��DT<��2��Ky��	F!�p�LxnϺ��U]s�~Ϝ���5��qv7m��FX-*���U�,��D��r-1��.�h3�w�vp�[���ݦ�yE������+���%F��hG�M5#sN�l9y��k�ׁ^M׮�S�aM^��fV|<#�CB�X�A��,���ߚ��#������q��Ҵ�k�f���U���\�7��y�Ӆx��ّ��b��E�I.49Y�^��뵷��uO��������c��@�Is&���=�H�,�>�K^���,��t;���J�1�C�#שMTHJ'��+ǯ1��i����I��q��[`�rzqw�^�5xvx.����/�7��|��jY�En��C����Ls��2f,�)�y�<Q�i���	t+���������u���*H�UWP��G�x����#�bO�5��u�T�)��T�=��!��Y>��H�工�i?��7$��n��M�Z����i_ЀwdK��pHn%��GYzJ�TJ\*L1?<� ��F}���ET.IZ��v�u:F�RYn$��U_l��Z?1�&n�Zz�f�v��b�����Sŭ��kKf��$IEu�S(M��-�܍��Y����|�tU@�Ĩ'����;�3A/}�ϩ�U&^D)����=@�q��sL_Kl��aP�kk��!f��=��ct��;j򞈢���^����Z�/^��έ�<�0��:�Ѣ�b��t .�
!���ف�2�c��A�sܠ���=�>6%c�6���4�?�I�%�t���J��dZƿ-�V�W[A�}��I1�6�X��S6Ѝ���Xm�
>3[�(�X�؈�o�м�hQǫ_jȪ}S}W�7�-���b�(;���<q�5�O��X��f �!$6E�Q�=�%�8Rf!��π8�h�6�Sa���D
�a^a͠�*z�Z� W
.r�¥����I�C��K����t���w�<�jt�l�Oؗ�`<I#�>IW��d����7�U�B�eJ��ݽ��~>W��8ݦc�o��w|'ߋ�el����;*x�n�H�s�ʖ��R[;V$c$-oOe����TZ�����G͌��*L�<8� �Z�ΡTyC�U�~V7�Umg��T�S�P�ڎ��=�r�!ʺ��m�<�h0�?lf�@�:o����Gg��_��Y�FCā�b����t83�O�|�|�V����|-����iX��P�������¿49��0��(�B�)�Ek�I�՟u%(��,˃o�Yc8!�sW��#6m�15:X�yN�����u8o�
H	���`�&��'�q�J@j��۰�e2=�6��4���(�E�m��jL�7��:��\r�R:/=G��./4+��"��kל��������� �T$QX'���Ѳ!�\'�Z�n�+]H_�l��b����J���0*B��s�����aDd�!�e���f��EqK�xO]�/R1|o�|n8mΪ-"ȅ���}7Ir%/�S*��Y��vnF���Am�sl���Y�x�u�N�w�e{N�@=7G�>�\�1��6��^����b�c��S`��Yl/]T���	�5(�/J��	��䂗�j�������{f�ґ�� K]k�@�jX3�>��������E����vT�O�<p�ge�hUe�\�ŶӚ���nQ����عZő��Xf�A��o5��.r�G�Dc5ց /q���-J+y��5�������� ���iIh`��bH��^No|���W_<7��Ղ�~vC�#RӐ���!tdR���&F��Ҫon�6IK]@�e�4�v����IVQ��(�����uH�!Q�O���	㘂y�pE)�m��QV�F��kP�G�\c�ҩ��S�ɈQ�q�g��u�O'�a��$�{�lD��>H3h�[�Aq�
Q��6�qj����cm��c���^����3,�¯����撊�]Z���!9��Zt ��`��hw5�b�D����jT=����N٬��ڠ����Q�4j�DB?���u�b��uT��) E�
Ik`���`b���9�J�X�79�"H{J?3o�tw�x��MOMl�FF��z�w��ip�`=���t���x7���\����k�&Nj�Τ�>w�i����W"��v�O)<��j�
T�����P�;r3Lu?��A��v���Vb\0���>5,aB��,h'�}�l�`�
�F=fed�T�3�釮������{3>�M�6�W����3�F�V矟�)l�$��X�(��d'�_`5:�C��5	�V2�M(,�LO%P�~��5�~¡��C9�a����"��@���V3,
R����!.������[�5a�/����I}6ҪI��F�b^����"�`�����������7�Ҍ�+�E�8�0y~A+��2��ut��R-����YN��`�/~�~�_{+�e�TN'�U&Ծ�
�S�0	����$p�ع��U�_����pH]_n3��� �!���F��`m�EA�_�U`ɏ/,:�h���3���y��׆B�W����|�]ZfH�0i"gࡉ7�d����̦������Iu�DY�+0l����j�����ɍ�V�֝�U�E^�M
n��v�
�1�V��������>$�p��Ǭ�mt�X�"��+�O�����*��ԉ ;�܆�7)�A��F1�Չ�}��JS.#�QEV��}6%=�PP�_�9���B���xʏ�H��� ��#z�@�
��\w.���w�Qrb1��=\�
�`7��-�b�C2q����n�nI��W#5uCvq�+r��Z�|S���2�$�]
ðh$��5ŭ����j%�&_]����7�����N��Q�8�� -g � �Eˏ����lٚ"X�� 6P�;�薎�Jߖ��$�G�]c���1�������/�a����P���]�Y3��<����ȷ�:t��g�JXT�A���*Χ�ؚ0��皠�ɠj���9Y�ϭ����%���>خ-�x8�����w��u
����A��nh��dM��B"��Ȭ��Տ~���HhC�Ժ�	l]D�i���,%t_+��E�/���&�_��0�5O�D���!����t��;snB�O���Ç@K��y�h4;�I�O\�5��Z:W]�a�xd��L�[���Hr�G|���(o�\���u^}�z(���n��n��vvH���&�e���E��#ph>���:�9�e�T`�c`;r�юqޞ�`>(	{h�f�y��x��k�N��?@r
�@\=HA	4=�|/ҧ�~�z�_�Ml��F�?<�.���1�V�~�æ 뻂p-�h��F��?AN8U!��h~�� ��ᓯ?�Oc�RP�r�{��:�ҟ�n�9�l D����d�������
�;9Ϥ&�i�pk�FaT����D��ߴ�JRN4�Gl�]lq /���Xyn�%�;j9e(B��ƒI�e]�b����c�@t#7#���y3�� ���f�V)�7�ȱ�3�R��38��$�t��D�^?R),�:�:}�Ʃ�|�?m�ܪ����U>ʃ��{P�ݼ����^�h�SHn �8	u"�9^Y*	\����G�N�_��퉨`�IM�;�P���2�*��$ΪZ׬'���y�f�f�߆�F��0[��Օ|s�$f=��_N�%c|��������#j/Ӈ�������u��h�.����z�ܜ���mLH101�7Tz������%�*��J7/�B�������q�N5e�p�)��1�<��eٶI�#�+���n�c�ui��wo3�~�ە����Y��q��i�͝7�i�X�u|����ف��>Uz�lz�ӂ7�L���ؚ��8u�O����'�0��fx�h�K����Oxh��20�6����rSI Vf�iL"���������=���7s��������k_`~�B��)\T��XyՒ?$��7����4r�?l��o̘f��r<���D�ަ4]ǜ=~"���1�-�p�ҞiN�B����î���i�ˁ��}g�u��:m\���Qn�w�k���*jۃ������(9�-)"�6���Qеh��9M����9;��t�yt`��x�d��t�n��.�}g�r?˺��َ'����tk���j�8옳� ��G! �o7KW5�m@k���T0x{����c�&ԣ l��a��g��A&ל��7 ��$�4.�׺����g%22�\�T)j`���9F��'�{�m���*!_u����|�lK�S�,	�J\S�KT� �Xq*��QO��#o�� |�<ӉY����ю��Q�s:b8��dr��L��B�!@$�M8-k%f��vJ�;:$��Uz�4<�ѽ-�F����<F���I,�:��O��⇌��
�lZ%�S�O��2L��c s�B�� ̸�C㨳�E�#�L�)[C�3K�4:��Wh��`����ƚ��m8S؀�!T1�fV}�N�&qo��ny�I>qN�Q�P�#?�+Ѱ��>����nVOt��%��V�G��TV�My�_��ȏ��O.�Ӌ=�7��n#����Z�'L�u�+�u��ny#�R%<?ͮ\(�P��<O@�D�S�c�Q�T]�)�,��-V����r'�^.&�A����!��E���hf�.�}���
�7.��C��vv�(1m%� Ι�X %]f̉F��Yvnk!I�v�sp���:����4{�觿�^�N/A�_,��ͱ�9�ٞ��᭚�*0�;�#�*��Lu7'_���=�SR��!��{��.���^�s팂�Kh����;��)-�����'݃։hh��3t�S M��(�lOZA(gh�ؼp(�Z�r��7����F�aYg[}ń ���	
�u�靡��*_/��eb)@f�ӭ��m�����O���7�|>��)�]����)g_L��2-pw5A�t�;xd.g�6 y�(͕�A��{�{�i���4-��l���h~�9�D��߇�n����$����Qt������B�W�S�{�h7p�^�T����&�`hh�M%��	މR,��P�)ɒ���q�u��̆��GG_��n$Ր˔�M��;E��m��1�L�;l�}�󥈍޴v��
z���s�?��F#�3!�a� "	qS���4��{�}�4)(G��/��*g����e�տ"���_ׄ�w�����p����A��3�̞ќ_���y�@��[�T}<�>5�/�����
��P��4��mm��A�e"��Yrֻ�r�I?�c�Ng1A�J����B�&�vOs,�˃P�;�s[g���^�����Q�W��|�d����Z�v#��3=�N��A]>Bpc{S���@�p�H	��8�� ����p^{{��JC__U[㇧b��V��lg=�S"�`�U��>�a�'֏�0��u����Z����,��ta��#�薱��Nw�f?���m %�lOH5�Mlj���\�!_XEe:�D.V� �ߧ�����2�w�9��R�����"���]�BU+%���y�ꆹ\����Z����qy~��#�2at�� N�K+����q�� �UQ~j�� �V񈌖TZ��<��E�_n.��P�5�\�9*Xfi��3e2RK(u{��9�?�@MH	�Eщy�{����/������xC*�5~��}�j��s�9t����e6��Г�+������M�#�ݍ=����Q���{�C5�W�l���C��q���4yI���{�(ܰ(�G�P��^����|c�Gb4�Ԝ���Sѕ"��������5e�W��'ޅ�����a��w����N�O�GwZx�lV�|T2�E���/���qB���S����Y۱��[0��vS�H~6 ��9�)(UɎ�T�<V��+q
\AW������3���m��p4���n|U�qB�܁�`�2�Ԓ�'H;�9?O��쉎�]�N��8[u$\႔�v���Vl³L[-�g�|B��'Xw�s�$�����NQ̅}h(�Ty�B��&�\u*�Thw�C�ZE� ��^N�7��i�r%G�	ֺZ$��=��C�Y����n,(u쿿mR�ʙ��s�)c�<�>�w׃S�@�ڃ!#r�_J�7,z�Y�`�BO,TνD��£��W�A�FgNAl����)la BP��-�w�2/O�j!O�)�o>\��M�f�{#�CV��+k��XBQ���������b�*����0$c��p��|C�\ဂC���|�q�1}����ζ�IX_��7�ݓR;�SVoT�H�F�iF�9��Ȝw���Q��'4�
 �x��*�.��5�p�D�,�E�c#������;0"Ec��s�c�ՏSH�	��8�]r�H���R=��n��DW���L���
��RP���f�Rf8�0A�^�(5�
���L+�]��T,e��O�� 6MJ-�皜���Yݩ�=#`���uf/�H�/�V���^�T�b�7cJ�p� D�<:�{��-�8|2|��6�n���=`S5Gn� �?�;�O�<�����1���69�Lޞ�f��6��-�R����������CZ�ԇ2kǔ9GK�?v;�-�@���~�7 z��`�6a�ߔzi��U͂��j�b�E�HiW��@�Tt�������~cPac}���?Wc��w��Rj\(�����l�jo;��%�?�{0*�Qe��Z�X���NReF����2�{0�5	h���
?5R��T���' ��N�/ݗ&�DU�b�.�u�n��w����5��ccevC!�����e���2�x,!vJ��2,�R�J߬�NPq	�a�#��m� �B��ڒ>�y�#��Ѽ�,�n��Qg�S���^��&^��~��9�F��$ׁ���]�*�!�.a�Abe�.)����:L��NG���`�l�����ea���̄/�t�Pc�S호~>?��0V���Ǩs�mZ��F����%�fl	)�k$�hpb�l�Wʠ����xD-%�L��ه���4�~�/�T�v�s%O���3֍��dY$ڜ1�c�ߡ�x.��i�0�?JF����zQE�}�4o�;e2�k�hs�,�N���Ը}z`8-�О2l�\A+�����1�*0v�k�%�Žm�)>�5C�=ƌ�5	B�e���4/,����yցL��8��!E��������X�=_�2H�dכIpX����f/���T��e&����tfGNFQAEC��U%�[����G�z�y=O־�$��{����N4@%,�)��b[V�m=� '�j˙\@�V] �]Ʒ��:Y9�B[t,&��!�����C&���Y���S
��	t�F�ݰM'����ktG"���m��i�+���dd0�x��:ɰa�;~E�C��{Rm<�*-�l�A�T2��=L4�q'�V�ж��5�8���-��fr/�H�����N>�!_����wѭ����6���^5	dx��F�Bl�J���W��Z��ycYw�B!��&�ۜ��G�(E�=����@���f��'�Ҽd�I�״�������꼄Rt&ԟY�	#H�� j����zIj.��e���㹵���A�!��(V\�x-�������&lg�F/f�)�U��?S(z΀ߍ�#\,���i���s]_�$��w�� #
��É���yjM6�����A7[�iG#���Vk�|9�����wv ���>U^2ٍo��i#~S�4A�� ��j㋻�UKr����4����QNYw�>��� ������+<`�3��GN����?��"��P�W�5\iςU=�&�C\G�.�
T� ��c���^���t��]��������ay��S���� ����HJJ�(��b2W6za>��3��~�Z����_��a�#�&z{T�~������K� �>�#��=�H��4����1<O�r^c@�/�d���e5��<�d�G�̋�2��I�u}�8�rΤ�g-�Ff�I~ؓ�h��!���b��]&��lY�_3�niE���b� �j�_�uî�u�jkx��a�P옩-Fk�On�:�0ߟ��p�i�%N���e?F�-�X�2eF]BO�2�[�]�%�2
����}`O��HHက�d;|b�E�9 =H�2��9�-^E����Q��y������7���$ᆌU�̝�Х�;s�fV9�e��1�#o�iؤY�}<�
������?cJR���M�1-�t�Rj��/z��CHp�?�$�=l������5�M���xY7����.`��S�፩"�ߟ�E�-����:�C�ߊO�R� �B	��ޟ2�����{�Ew`�"�a[߆��ϡ+/�wp���_�ڒ��e������7��N �j��8��.ay�d����橆N�2��z�aMvi6�;X���Km�3���Dk��ZH��� �����5kK�P[�YbԸ���������#ͭ��h�C|����*�5mE{��d�Ho�=+IB0�3���IG݄�D>�W���#&�|Y!��h�E���h���C��j�l��Lΐ����`��j�	{�f�g;Ew�㨤�TG>�����b�b�����
'��V)���I��A,����k��d���U<��L�	��6�c@֧)e ��h���?�=�����tp/m��N�� -�Ep�'�;����j��8�%�׎A�{���{;���[�Ui=4B#�W����qʅ0��o�7\MV�����[OO;pAz��0D<ry"0���`�|j�*�p~;��N�j�[�
M������k�W��/8�����b�\mrZ���l������K�i�(��,�DS��K�eD�l14����*F�3A�?�O�������0֘�_b�h}�p��A����n���!���1��B��'���5�O�s��8�@Eu�Nv�j�k��B{��ZY-a���=�;�(�`��Y&37�F�n����=̻�i���p߅��B���{� ��z��zD��c����*��y<l�#��ܨ�� �]�rQU��m� ��~�IMв]Nrw��Ų�q���d�O��� �6'�Fy������x�_�X�]�D��U�φ `�,s��7��: �VN�[�@��t�T׾Rz��o��#q�����8"v��.P�B���.P<z(�	�+���͟���d�q��,���4��?�qv�X�k�hK@H?J�>��O�V{��V�2:�iB)����	D�zеvi�/�p�4�;y�a�Ԃp( �ѵf�o�y*�$+����Ѳz�!�,�?3LZk��-�T�����)�A��ޓ�xf�/��u��VMQ"��+��V�^�h
O-}������7�&>T�D��+����OJ�dB��B�x��-�E�!!���o�f���)���A#4}o���[e�
�����f���ـ�&��F���O:��`�mO���d)産�S�-�0,G�)��b�0^�� �=h�^�g�:|��ӆ�y���O�#�1�
�̈����wa���6��Ч��,�a'�w�u�$��2!7�����]�m��u���������_�$z�+1�� �Q��Uv-�z����a�N|��V����%��Qy�`Dǃ�!�B�!]��&	|��&�HgלO<=��q2��W�Io�.���K:�E�^޽<p2<b#�x�-�B�`=�O���^8gWՓ�嚽����~0��3�M�������	�c}57��`X�:�ثP2��L��2,K����\�Y�ˑ�ME�0}.8�#��+$jB<����Ee�5SG���	k����vi�����\P� oA��2�8v/a�՗�U��(��q�5߷4	�SO�&Dd�J���*����N�l+����]���+����(�rQ� ߧ�@�!��P��.w�J殇l<���׀��$��Nr9JKgM*aKi�}�S�g�)C(,X~"W�u�Ml"��S�<��xettXYQ���¾��\�搹��̠F|��\� 6���Y�Z����N�����KK�c��>���N�\HX�0:�X=����6��	��D~"A�q�-�yeʀ�����'����UO�
�v6�T�j�>�����.:��T���Z�9�ц�����(BLD��M�g[cGZE�+wg��Էz���e�u+����/(������"�^):b�?��R���1�IQ��}�A��gbw��%�/q!���a�<;����/y��ͨ����Gc��)���&[��� ֕�
�iN�� ���0!���椢�ZJa��}�T���0$M.��ë𘏵���DŬ���:�/�
/���s�����|����yU��3��� '��үzh�d!e��^qyp�D����S�|"�5������w,)����7��&�)�n@6���47�E�iwҘ��Ոr�Яn����#������F�`Z��z�Ѱצ�;�JR丯1>q[P�L^B~���4��l���vB#;�P�pi���C�~�j>n��������2cީ��xv"�3��EN�g�����n9���c����MA&��&cG��>��3,b(��Y�w�#h����9d�M-�#I7����siF�N���� LO�8Tw*�\e�n���S@]\y��u�L����e �����R@�����jF��fO���W���0�My�Z����8�R�/Sx}�п���Mt��VZm^�����Y%4���?�b.0mlR��v��f�m֚�`�:�%����"�<�^p8}���+��c��/iu�M�e�Ռ��z	��f�`�� ���+$pz��U�\�%�rw{��W�Re}Z:��8��Z�~�G>�]]�ӈ�i+cc�������\��͑6*T�~&�V�{^�}��(,e�e¡����~�Ο����+�<w�����tQ�6�:
ޠؑ웮�c��i&VrNDAF)�/C�uTc-�]GK��c��:��0YhnDd���D�!��B�j����C��f���|��W�͞�9��]O��r��`�W���`j1VF������'��M�M(i�ŀ�KBX/3��`5�Aw3�<��J��P:UOP:���4X�*,� I��#��{�{)=�,�
���>����a���s;o3�o�Rѩ	Y�(�ZƆ��L�U܇o��B�B4!����a�~�
D����x�܍�B��2�����+;��W���ؔ��粖����ˮR�V5u�3���"x���� �2[H����H�(Ȱ��[K�)md:�^��h���Ȇ�5��������ٝ�N��5W��t��ʄ?ٸ�䉍�v��x2�L��MZ��Od�&K�R��<:�W�y�9�����j�׌Τ��̃=.�xY�������%L*�X� �/�3������ꤖ]k������?����W�Kb��|�1�[j�v�	�}�f��^��M^÷dd>\ �-{�ׅ��WC�4��?O��kޝ j�n��ٻ7�=9��U#���3��7���>r��1 ߑ�Ӷ�Q��*��^.*���f@��0}JHg�Ng���,RlMj��j�����j���TB^#��c��i��x���0��v\H���z��5��f��r�EJ��H��z���A�)�=Y@��P�� �_��yH;yq��%|ᮝ�i����AO����᎕�D02-�\��I�������0�70M����*l�]����뫄���D�;����>�
�?�v"�q,��.��M��
3�����8(-AT�p��L���U�Fq&��3�v���Ö#d�L���)���	@�H"O���h.Kr��
o3�0p����(̢R�[�fe��:�)�ջ�>B+x�R�s�'���*�Z���E:5I[8�����Z��^W�k�^�<��b���_���
	����6*n��N���a��;9�{��,���}*�*r�	 "2�nչq����M�~�)ؖV��F�7�CQ�a�N@t�����c��;�����B�Q�%W���]��� &���h�Մ!�=f�	�\9R��!�D �sel�����]��]b̙_��ͧ���Yq�w��MY=�D�����^;~���i����q�3
���	�*Qi(�Sk˿�H�&�N�F)[��Uytl�_�Aq_X7�vc�6���վ�Ef�ͥkN�M��E�t�� jX������wW���t����̳�H�Lo�T܌���dй��.пq�u�9���,�V��� n���<���%�UP5`��z�6FIaω�#t�]-�(g6�W��w��2�h�����b���؀�p�q��z�̦�2�P4�Y��"�L�������w�`[��N����		��iVt��C��u0����6 ��5P��:�@=����W���33lo!����{��V���UO1b��W�@��ro��j�c;�ͷZg�Q�<Rءq��(OO�{[(CA��V� �K+��,���5�K��OV�@S]W�M<�B�'_�Y��g�=Fߍ��2:�cĎ�#ty�ͧ7te���w����L���:3�%����L�a}f"�`�n:6ngW\�����c9ڽI0ܵGR�7)��/�;Y- %��x��V"1�c~45 �����0>�-�y�Y�ygH������l��9�P٫���1�^�@ݳ_]��|hZ����:�/r��'��pza���@L����w~V���qr��udU���	d)�!M�F{����%�I0�;�8�P�������o`�ضmJ~md�%�r0R�~lc�����>�=�Z��5" ;	m���w�pA��������E͟���~��/�B���l�1Zr�L�욉CAb���:z�G?L\6IC�7򈣁��:)`[��O�m�O�̩���?��ps?zN�̺��DL��W����~4�k4���Z3 ���lY�}3\��-q��;�C�ճ�a�ոFc��O[!�%�]:����\��Esh���!9�DB_Xb\8`1(���E:����s=��B�����ط�H�G�&B��t�N�4�ե��@e�Gy�ذ����3���Zkk)�u�gi켲��,��Eh�a��z�
��֫��!��eIT�[(�in�3|��7?,�4�`5L߬�݊r����熲���Эw��	��w ���2���&ren�#v���q$�x��ol����y^���j�r%2��&�] uc�ߌi9��yϜ�Rqu�5��nP�7����W�N46X�4k�Wpg��εZ�닃���&*�}g#���U)�������pxQ� %R:�bClqE���m�O��',lT��v���to8��]AY�AD�FZ��+�v-w����NG��>�D^`#8�2I��a�o>Q�wP��YDʟ�ea�
�9$���β�G��������>�
A����[�TZBoE�S�`5o�T��e�Q7t�o�ovO���w�ѷ$7�+a�����?��b�T� �a�7<���bp�NNe3�ظi*"�~A���z�4�xxH���7��t��#&���EE|~"`���ԡ]Z��$y������*p8(Ur8^�UB�����?���P���m���������d��{�R ���eda����S'�rc����H���I�|�Ң�_�N����\��F�G�t�I���T�BP(JI7r;y
���ix���_���8c�;o�$�ro$�喵�ȷo����ڬ�H�UH1!���S�z='�3�җD�؋���!j#���6%a�!_'�W?nL+���չvl�/S�B�8�M![���9���A|�DX*k�+ ֵ��&Ԗ<pf�*�׹e�類,<pI`Rn0����H�����t4�J�6���d0d����\�ܽ�fo½��p�E���;�P'�0��&�����q+�p�5B��^E��K�a�>Q حAy/��y�(Ć�Rc��Er!70y�N�����Tk��19�(�P���5�AY���&�$�����rj��a�� �+�?z�3ԋ��X�4.�h���i�+�/�0�䋶��Ʈi��.���DiZpS��<� �e7��oR4N{���ُ
��.�M)�πr	.���0�� 6K�@�iP&�����4TP8���PB\~��ÓE���KP۪ц��ڳ��-�m?�E ��wsB��k�@�dk�B�=��˪p�w\"m�<j8&����*�cv���g�|\\���%z2H���<,;r�[��"��4jd�(�~����E��Zq)�l���㍗�WM/N���,�r�ڸ�$X��?�ŹK�Q��+�u{!w@E�}_ŗԸ�a��i��ОW0ͦ(�>Xva\ơ(�>����J���Im��l�2=L1}Em" qQE���HV*~4���[㯼H�5�ni�8R�:��U�����7��{�~����w!_I*f���;@�H�{��e|���K�k������V�6T(S��sJ-�K�2�DK���G�{��v�`�۬
C�<�����Myz�X7���rM]ߡ<lF)��h��<��;َ*�n�Ν�J��U/��d^b�Z9@�#3�cx��~]ͲU��+Xr�]���'m��~�Q�r��;��mh ��i�,p�a�D�^8Ђ��9N��è����Em�!�Y,�G=�8���N>��*���M��ב�\��҂#�]�8.����0N̯�Y���/�A0�?⨩�����#p���ؚ�#3C
#���d�g�5���]�ޅ���O��\�)]JO�����= ?�l�-��k,�h�(�hlY�&�3^�8ĉZ.� ���-*ʵ��0�s�S��+
�'Lԟ�]�vh�uI*�흅� 9�;>���I����� 
��"|6�C��qD�E�B�]0�Q�8���C�֘?|qtd��-����������9xܺ����,qvi��A��wA����o|L� ������p
�s�u�H莿��L�1�A��\t�%R�t ���+ɏ�8�FQ���S84Vt(��#O$�;�ޘ��N���l������~6�!E�Щ����s��w�X/�ڽ����G��V���V�x����H;��W���r�.�m+CN�RZ���<���4�WkS̛*���w*Hh�ؠ�tq�`C��i���IE;%�RA<u	��Jx�g��6�y�!y�� f�����Ua�(h����9:I�η��f=��/>JW�Z��9#�
����_�ׇ)����^n�ߞD�J����ǿ�,����O��t�"�˕�P���ml��/�������9dw�!���D�^���<YXW���ĺ�53t���&|�Mm�g5�������-��$wi����-#���l��������x>�P�'/���qq�!�����5�j,���E�>��w���md�S��s��j�Y��N�+6���1ڷqN��U��Tgg�������!ߚ:T�)��nx��t*���~�[	=U��bI�	�b��)S�Hw-�U�J�M:��*�j�3|qO�f��t���,�#!�'|�oo�Wz?���Q��}1k�!�E�^O�z�����m�k��sО�n�2uZ7���*wL3~h�?XK�ӈ�!Ro�kNul&4W�"̡\�+�u�S���d@�}�%~�3!3���{K�I|H��}��/�<�θ��ư��f�|c���U�s�)���)��54y���u��?O�����Si	���aa$�;�}�W�ρ�#�f"��|�Ɯ��(0��?�# ��iH�[ ��M0`��%ݝ���'�d�^�Y�z��K�EZ/9��OQC������L��fX
`Q���@�@֥����E����b��<Vs�Tk�F��_0�d�4,�����C�uQ�H���V�㊏Y���~�k@�[�ȸ���څ�g^��Y42��GV[�M�	h=�ιJ�8��f��t��rڙ��N7x
[Ie��\�, �v�T��N;�Iҕ�lG�s͇%��?}(;N��rBh�L���3�` �CllU-�+/��w���xC/�������M\���\��n����Ӿ�(>�u��?����U@�O��q�h�"��'v�c��3�mKo�� ��5�����7[(Ĭ3���^&/����do�߯�#���\3Zhg����m��NciL�>����.Da�F7��?�Wrau�:;�;'L8�'���t��XA��h#و����Z��S/����l�J�?^N¢��[y���� ��P�@#ߐ^�P�ß�zq���	�A�c���H^�$��`�v9��7��,eSs�]K*���W�V�ސ�)l�`�+��@�/�	6��u��Ƅ��22U��[{�%���jaV?m7���9ȏ&��H!�� ���,��k�+�j9/�N4M��F�݅��*���7.�P3#���W+�cxF��!d�+�;�쥋΃�ATO�R`�M�,��.^�JY�~a�2�f�U�	�l�A`�� �����ʹ/��XW�?s�4�&����ԝa{�"��;[l��]_�����%C|�U�2�sj�9�tb�e_� �.�J�A+V��nJ��j�b���e� ��5�
��m%�v4�|�����]��z������6��	\&��lU	M\�r�K�Z��j����Y�wln����e����u����On���b,�`��6�f!@�����o%���A܊`��^u^�-'�o�`����D����A�x�o�C�
o��
���$����.`sT�{��i��s��B�n~qx�AOvMy�̿.���}��e����}��a��[�gx2@!�";�&ա��'9{xɪ-f�Y�0FDg�vd�����K��(�(y�on�E�_E��-��[���!&7k����1@8ٕ�4��u�m �dG�y��u������߰������YG�=�r�e�$",��-^��]8�/���j	���&�k�}f��I�1��蛠C��q$L�怡G=�쫆�tP��6�z�{U�>��1 ��9�V�B(TN9�ʼH�<a1���J� ���S3�'�lL�kO+%��G0]��M˴���y�CJ���:�U�,�Tk���]^ � 8y_��i��wڒN,D��w�Ϯ�W�?�|�ʓx�l�����d`�VD$IY9
�,{�i$d	@�Da�yʉ�J,��ĳ��E���}�Jk��Nn�sH�s�����`�7a+9&H�D5��۹{�L:/�Q�w�� ��P�""�(b
K��q}^LӦ�����w*����!�5iu��v�<�sj8z����#8��JYׇ��e�����+9EĦ���HHm��2�
�2��Btȅ��Sd`Ng��t����1q������*�6�ij%蒓���<a���}ZXf6�"|��X$����0����z5�X!�_�U7X�^�<�ɳE?�͛*R�X��s��>{BM����yA��3��x+�Yŗ?�iχ��k܀�������䤝O)	��$7v\©,��ț�dW�q���Ű	�
��U ��{��>֧$�猬_��G�#,������Cv���q~�a�IM�d�,ڡgCX��QQ�<<�P�9\�E�:w�Ms�8�z�>mqDy�S6h���$	���PwH�'Z��c`|�y��O<�0Y�
��5��ki-2"$0)�ʥ�J�
C�du�O:`�:
ܭ���;��F}���������T��q�;����T2�y #�L��(U3�UF���)&@�Pf�䔇�KV�N.۽�+�W�E���ؽ�@�E^o���j|�m��b�qW��䊫�|*�:��P��8���8[��Ǥ�BW��<(oB��X�߷%�8��|s}�즶T;|ٙ4)�����k�S�O���H眮B�qdkZ��԰NR>���X����j>6ŵ@��#;��P쯜�8����X���x%_����u�w!2�G{�ޔ��A\r0
P܌�ay�]��LM�JV�\Ե�H����wJ��ꋎ_7�%�
(\
deb�p� B
zG#[�,(�%���Gv�}6��o:n;ǫ�4)oAg6��̀|��(h�_O���d!\�T�Q��2ߓD�~�(���#���g1_�'c�2B�k�,m+�����M���wS9��րVgEW:ߤĳZ�)���Ħ��1����M��g;�\�0��ǭ(�u=+$i�B�z5$%?��Nx�o	��I���E���J,1��P�F��[-��k��D*x#�Kυħ�-o�|MA~��S��ai�>$:&:�|�X��@Â���h��`����Y9�=�}]@u%?��g��v߾�uƣ��(q}ዎ6�L��+����U��
4�k�H�?0H�b��0���k� �ʎ��|�� �����9 ����u����Q���|M��"kD������t������1�%q{-�� G�4U
e3��¶\��(r��@��\�Z�D������Q5�I%�Xq�!�I�.��w�,S�y��33@�RF�3Ӛ������kf�L�H����̓�{��p�����<A_�;��@����2�wEh�O�ih�r��> $�]�y��L�*�� ֛]I���d���`y>�ĩ�>[�T�چd���؂o�/�/���3���o=ee�o}(����f[N���=W��y�?��?KGS�ؾ(0��"sB)�6VǼUm���L0��WJ�j����c��g/��?�S|�@�Sl��ew-0EG�m'����:ۘ�:��/���S�a��u�,OdaT�c����0�hX�P��p������۲�Еŧ�Be��c�T8�U����q1�|���?a*�b�H`s�Ou�l;a���-_�����M�d�ۼ���K6e�j"(s;��@��{dQ��</vxOS��C�lm��)L��6Ɍ\��&֬Y"�l;n�/
�_� "w���� sNWn{!A�9���~`Hc5��b�c1���l*��"�m����������ӡ��� � V��ق��K�@G�Ŏ>I܌�j��p��%�B�(���f.�*E6$�|Uu���T�|�`��T��t�����ׯ�#���T�ܫn���WP�zj���]#��#(2~|�ɣo�[���P�o�zLq�A߄�h�@Պb��2�MI-a�B����G9��v��|%�v"��a����ݔ-���$�dr�Bm~�>�R��΀{/��uG��L[�Bp���6�}�FS!�O����ݶnDzO���n�����&l��֍�����Hm����/��#�Ң6!��N �8�Yd'�?t���ή5�y�Z���w����m��:��Y�^�v�z�nttTR�����{�����f�7�~�(�70칹��.�Ѓr��s����>`�͓��T��Razb )���8+{ݽ~.K�|�S�&�t�&�j�?�7�nUY�]/vg+E'�ś��	,�{�Ƃ2�qII���'^��Q��=�䌖�8N�(�>�Qo����O�X;�~\<f�
 \����N�݉�\Y3���T���^����>9�?�XB�;>���:�E��kY����@�D���~���lL#*��5p���	�̇�g�T�H�7?�)e<7�?/Y�h��m�¿��Gݍr!mt�Oc�N��K���yeR�%Q��k�Mw��	!M��װ��Z�?���V���qe�f2;����)�1N#�1k����1RX���_8������O&ε*�,�ӳ�p�*�c6���k��Hd1>��H�?H{k[O��O����{���� re�<�r�4���X��m�o:hs�M6R����;ꍙ䨩\}戡$�ӈ��z�A!/\�ǘ�_�cЁ�7��Z�3��l�~�S�v]�	�Y㏛�p����	�X�!,��d0q�"20z��f��l�L3��a���]	��o�&s�)C�+�ސ���w���h�&<O�L��J[{d�kX9�5�=WMnZ����ǀ��ER��)i"B�HT^��u��?�:��VT���h���@]�D�/`��dIl�y�[z�2����p�{��Q��8�P�m&83/�J8MV?�-d�����F�F���{[�BEt��b�H��L������C5�]8���=�wǗA"�y�7�b�����Ю�i��*m�Sj�F����qaqE�;mq6�'e9 k1��D��g�k���m��-�����6���Xu�t�c��S<��?�)�&S��I��_ FZځ�
o+P���EXQ������.��q��s%��E�F*7=b�YYr��HzQ���s��j8�]��P@%��FC¢p�����{D�^�Sy{9lޑub�6��T��e�\��:�˰r�����R��u�i�/J�2�&��*zxQ\�+��ԭܜC"��W�;4�u�I�c��^F�Ӟ�KP�{P�(�,�}�����'���Ƌ٥�DH0v�i�>3*ɶ%�C`J��Χ�s�d��d�qɭ���k�� �b���$z�J�[�e#����x�<c+JU���Zy섅Q80,����OxS��=(�`3��O���+C�ꉗ[� ��:Y���moK�m�@�v �Gi�E �̜�ݗ��\�=��=��BgD��߽`�����B��*��S pS\V��ʲ\�%:�m|��E�*9�ٯ3+���qf'j�wSsF��f���n&K�w�q ��K@�nڏ�~ P[]΃{�Y,�헬��Ӆy{w"��K�~���K�Vi��j���Li��J��J�Ž��%HK�BXa�,�b?'������ﻴ�؅�1g�v.��t���E�tG�Q	:Z ��?}�J�����I-?����hT�
�l�F�ő�J�/F���0O�R�G1���-����Eo��Q3^$��E֫�:���49�fl}Z(�q~������H�MR|	�Zp��<j�wr�^�L.���EL���@���!� ��Ŋ}��U�m�<����X�Ί��p1�[.S���~����(�!&Ž�]Ԋ�aT��~�Y��t�����v[�[tq�=B���H]|5
�Ժ��HOE�s�/fk	L񩤺�+�L7P�1s@qscD~t����H�5�X��Pz�K5K�X�ڇ�[�L�q؃uγ�QO������^��[�
<��-ԓ�4�!3m��i��S�j7��IsTqni�����s�����
��\xm������
1�*9a-!�\� "��0.S�OF���Ip	�mCn6E��,q�1l�v��b��^D�fm]�l��K�&���L�)�!���~<�r�1%ةX|�qj�+p�N�C���%+huؑ����h]�w�P�������,�ϚA�M�`˷�p�0�rA��u?�!)i>Iu�r9�~�01Xش�j5E���
�SZ$�_����'�LQ���R�����æ�����Y:N2�<<����d8i�l��:j3�*����*�d�L��t̲uT��q��]\CF:bb����?�v?��n�OF;���/P�S/�kz�8�K�����*��ŨE�G�9b�l�~��QPs!���p�v�@��Փ!L�t3%h,_��K�3L�-op`��"��JS+rnN�C@�Y��Bnb !��>.{���|��
T�۞�O��U	v௹�R�x��<��b�*n5��<����<����q:Z�������ќR 0��I�f�D.�8�
MP� а��l�<���|8&�#�B%��J��jME��>�ID�8��	���o�}ѝ	��7b[��<3@�v�mU8�ZX����O�ǌ�V��4����{�x�
���q�	/�o�].��>%ǔR��W�P�qM^�/}�9_
�H8B*��c\%FԀ�0�t8|c#TB`��qNA���?�X�}˽�K�d��2�Y��;.#�
9o��t>釬�kYZ���e���&�����e�چ�C���y��,!���&�`��,7p�[U	�q3�� r�����?ڳ�ψ�9xal���a�<�?xܐ��U�=�<~��;�#X�|�V3פ�HM�.%V(���_2��������<��Yr�$^I��,Gߣ#x{E���!q�.�m��OL��U=����n,�e��dH�ׇ�H@d�T���J�Y��ht�V�ӄ�~��,23o��f����D�ǎ�6�{f�Ҍ}�@��@��=�-*)�e�L#��_�P[��,�LNۅ�h/��uXdZ��Gs�I�Ce28��qR��}&=�覷*��uc�K�� g��u���Z�q�@l`�8�%�ܢ���ӡ̆��D��W���E'�昼��ރ���g�ֈT]>G)���
~���������?,80M0?	�o}~�j��Yٓ�Q����U�����u��,|<}��՛WY!����Kfq���Y�{��)
��<)��OiB��c��ʼ�|a��D%\K����K�A�]�F�rȐ�����+��o��w2������zn!'H�:<�P���~�@ 3�m�r����#E���M��RI���m���(�ߊ���7Z��d[�������_��t�a�0�Y/�u��H�
���Z$"#S��ۚ߸ �{B��
܉p���m0BWW d�c�c�M�>$�ר����;��z��+��f�T�N��ALO&�ퟧ���'������k�<�]P&�"V�64X.��E��%T��*��{�{�jh�t�SK�G����7�#�(.�mz����j?����Ɗ/7�eP�¤
�O�3�۾��EzeA�^�^T?pؖc��ѻP)(���덩G�85&
/^����Dum'��HY�K��}�7�;6�.��\Y�p޿�|�6�m�o���k�&I �_Q$�0�6�i�<�!K�`�S��u����Z���2��-��?��q�������$�gʩ����E����/ͳLw�-቙ʂ��Y�
��|��#��}9�7=��Nh6N�#��s��\t�� '��P��ԗo$К�������{��<�m�h��a�M���00֛��+#�`_U����O���v��N ����� ���N`�\������Fh{0~ƃ�w$k=�di�N
ӧ8c�[���
k4F�T#�g&r&�¡��~�"��'�C��V�-9���ߣI=��8햀Xg���`�o�K��BՃ�U,?R١�6���\'ܿ�t�צX��Nu!��������^��ddh�Ly �q�������Q�׊b���,3�(����M^���x�s̩���J�pC�X�
���h��-q��)7�c	���x��]d������	"�Be*	{dov���tZ5qV����|�@b�rv��I�7�$o�<��h�#=cg�D5�ppyd����Y���Q��p�Y�4�p�2] .N!O��w�T����
����m΀X��J�ӹk�QJd��J�Yc�*g%Y\��i���eavcJý�EŃ�X�b+�<#��oc�n�c_�E�>�ʖ��,&W�{HZU�C
���G/f*� ',<.�tD,Ab,�]e�M�'��~�j���O�8�&�t�X\���.L]�����)t�d�bA��Ԧ>mKL[��B��2���ș�uO#�2Ɲ t�g��Lnm��DB������M&��S�TZ��h��#r�x��,>M�l�sp���~�{��-3�/d����qJ6�[|�gΦ����o]{�
��\��OC���ԛ����S�X�����wXI�� ��J�ar?H�;��l�Mq�1���,Ra$rA�Cf��� ��#u�R[�H�f��b�����p��׳��K�l.�"� 5H�=j�V�y /�7>%�#��m���0���R�ؤ�ws/���D<�H�Q	nY��r�~�%��qhj4�Ta�_}�[��І��1��z[�qS���4��\����[�*��V3�L9��4�@����5��l<�B�3�
�����I��#� ⭊�pM=�W�
��,&��Z��o��`��r>D?�:+U~�$P� t�o>��k�A;=��ׁM�B���]��k('��$�='��ق_B���	���p�oN�fT�
�[%���V��`���7�APJ�j�5��IA$l͓����@Kӿ�ieg�����[��?�$�=���#�3᧴xj����E!�w��bʳ�a��-Ou�H�n�%$M#9GT�ظ;M�:Ɉ_T쌩t����s�!2�#��Ӝ�c"1`Ĥ�����@Lp`��8,�����,PX�F�����cL����)f?<{'x��%�=��Y�u�����ci}K�d?�L�=]�"���'���x�m��~�zQX]��$
_�]���x$�ƒc��q�PZע�{̬rO =����ePzy;?���0/!5�Ձ;B�9t�w���Oe@.��
�`��p�p���MuҒ1���|!qkcr�P����k��T�=�8NX���������]�S w�h7]-���J��I�#��%K(�v����M�?�Cc2��:yN�gt��ա��nL_�'���1�eN!�|��H�}lp�) ���T�%s�	���ge��L���ۥ� U��YЉ��6��7�!)G��ݨ� j���i�S�I�Ӂ0J��� �3� ��l�	�p�u�LsX0�;��Y�cMf�O�g�U|ۋҾ��j�����w��u��iz�"�����ZH��s��q�p�j�����VV�c�,��D��AY�ɦJ�VC_�����E�$�]bg�D��L��cgB�r)���6sww��V-��F���wtE{���u}�[*�P������,R��H�R/��B�c+A�i��������@���\dY��bS����\g�� �6II*�Z0mAEb�Y�g��1���j�;m�E�L�����d�iy1���㰱��'�S�d�{�l�"���&Oq\6^�j'7Љh�a��O oO���E@'���tfqlS�7d`�zbǇId�����&$�I����b��p�wY��6�@i:�����x�o�R�y�M3�>&6� ���r\�������٩��ۗz{ґ����/޲~\��+P鳙e��BÝ�q��:�h4�~��z�vr��,��-���!F��.���`��A���ι߂Yv.��fЗ���� s�����c�0:F�@�XD��������TR��l4����)�t��*��[��1�����oSp$�M8g��ة�mS6�ci<��뻪���H�ד�$C�q�ݮ���ڒ$'��w���@�p��^�`S}&6I���p� ~�*��$~X&6$#���2kK&��yM]�lU�J>�0�D�R��N�H%�t�K�ң�
g VS��|�3�"����m?{k��\h��3�quaI�(����د��i4�?�KHQ���24ؕ���|�8��	�;�/�8Z�Ș��:�iV���#N�<�������!'[h��~�i�mC �XR��Z����K�k�W�$�|��.�toD�	=I�W���hG�P�:�o�����]&���v�TH�����:F�hvS^��&�&%���n\�0i#k� 4Y�n�T(b��r���m���G��(<���t�g&�pǝ �I�,&��C���	PX1�,s��~v}Ef�/d���ƙ��%�o >��^�>��-ɇ���a��̄��M处�e �����#�h����n-������ؿ}M*Цy��M\��mx��_�>�ƚ�T�*t��>X���� �o{X�>���4�^{ب�c��f<�^��U$�@�i�W��}�;b�������߭7ِ�@%��r�=���8��l\'�\,kD��ٙ�-�8W����%�1�y ?6kL�^���s@m�)���	=Oњ�ˬ]�r�W�@��t;M(z���k�V��o�{���lee,��P^��ϗR�
|��Po�@p&��v�	�`�B�k�1��E.�Jm������\1��N9{��7Y.F��1YȖy	{ݗ�!��=3U�|GK�X�܈s�����r,u���J��:H���M�O����v������UWy $�Uv�VH}�a�z^k�"��{��s)m��Y`�X`�iZd ��R6�m����G��'\�2�����bE8�юU���o�hdI'u�T�V\q��\8���Јb\ѐz/&Dd��/��D�
��l�Y�*��N�q�#����t���p�&.�j��������WT�꥘/+Ҭ1"� ����a��h�T�-�r<�8εe��D��U��]�{`p����|#�y�%����_r3�+��%L�t�|��uG3L��� �VK����y��GoS�U�>��ei)A���R�x R�O}bA��x̋�.Z��2�]��}�I�42�����K�h�����C%�F�e6��o��R���_\f�{���jB\�9��m$������?��k���99c�D����������f��$���a�n�
�W	�8�X�lj�|��/�c�!������/�J��.%�<����+@,���%�P�H��,��
��c��t7�I���2�V�m�D�WuT��[M��S�3d4R�Lx��]�s�����2dDhBx�|��u@5�2�| ��j�s=x�����2W��|��<�Կf��b� :�����]:ݦ��~��4i�VӼw���i"�̨��w� �67U���"�����8m���T��Oö՛G�V����J j�vs�
�!��4H�`��%����=���?�U�	"��N1�<D�ÍZ͆͸ug9d�PC�:�kw~�.�GFmt>��c��#��s�<{���z�k�$���:�H��[��
�HE�ۯ�';�,A���6T 34��[w����БB�Ԯ*��� ��R��K�x]���4�D$�U!p�f�!Y�>�0%:x�}�jgc}�K^"��X�튻�v3��������5��6Z�j���E��$��oA��˲X��P-�l֣Majإ�ͦw�6��5g��ԅ�h#�h`�7���P�|�%arRhM_걌��:#���ʚH�~;	rB	�am�Vt���A<���pN∆�����u>��GPa&��tB�\�|jO���y�H���^��tTm�X��ۀ���g	��e?��#<8�!��F����S�_���?��e2��T/֞(��K=�F�f�'(�g�N�
Ijv���*�b�֏;� ���rȈZ����U>m<&�=2%G�u0�U�wI���¶��t��١��e��=6.��m�d6 �_�(�7ݞ��%gkh���n�-&қ�?9��*�_ �Z��*,߮HT�*(��k�m,��[�uR�7#�7������n���'�!n� 6����Iۧ��P�X@b5_�c7u"�I�e��N�*�T2���f��砤
"uJ���y�y��"��@�<Rs1W��L؋��k��4;J0�	bg �s�2�[
>�iJ��&�6��(�� ��
˅�0��o����{�f���yEA�,a6���C���������f3�D�|�vgR
&�-�_}��Ʋ U4(�f���஘�����Q�����"������h�s��N�����R�z,U�����[+�Q�U(�)?1���)/z{}^e�r�t��y��Zh��QIcS$�gO
9z�T�*�U�-j��^��Kt)įwm՘M��^��\��z����n�s���-Gs�}�C��)��#R�/b�7�0�:�׎��Z��,�ۗ�Yd�Hi�!!t�H]�tɸ>�/uZ��i�q����X�7�Z�e1~�B���J��*���7B�W�$u!��_?�T��`��ix�s�����}<TB��:����L~~�J3��Q���Q�+�Z�w,k\������OW�I��Y6�a���ڻA��*h���'�E�m��ȥ�[7�_�I��u��U:��&��IL��I��P�@<����8[��?�گ��n�eG�9���9����n��V��gcۼ���N�n���Ѧ�B���(�u�1���iP4�)�|�q~^�`s	�X��l�g���E:Hg|��3<)��a!�a7���ßR�ݦIWau`x(|�L�b�z�{Fq��X��P�4K��3�o1�/�*�UD
b��5��o"<tH0U�_F�8�:,
j��3>�ȱ�5��F��@~Ni�|�o�g.<(>R<����@H�x��/�����1��*[�m�Ч�`iMYi
�np�:�r7X}�bK�Q(���%l�.���'R{����{�ؽ)nb��0�BB��F|^T�ڎ�w���1	P��<
��)_��I�w'�`��v��y�M#���Ҭ뎯�:�f���?��q�-�W�.�z���b0���	hѸ2f����P/�\��{�)
�}�"��S곙!A����T����A�n�կ�y�[Y��Ec/I��_�8�,��ĜDTS�9��L��=͞.?��= �H�Y�;k���	=����� ��/WT�ų�$��H��^>h95�`��xm�ѯ��+��.��-�H>��]�����U��x?�Q�>�ǁ� w���<<W� �r��`�ƙ(�0�˛�&t�R���[�cdqy�{��������JJ�9$��"a��n�mt������X< 0U �l���k�a�d��tO���SP�5��}/�aG��hj�sp���7�̖g\��U^�{'����+G��o.	L?�>��9���ygN������Òn���W.65>IxLzL�$r�&�i)*��b��${~�#�Tr/��������p'�bt�	P=f2����Ew?�%��"�V-c�U}�p?-��zȀ9BE��}]��>�Ӑ����Rh"�?�m��B��x��P�I�4(�}���Ĩ�(܏�y�fԧ���u�$��
�^��ʰ��g�� 8�� �HG�k歏`�8+�U���Ã��
@(�*-�*�+�����9|��Fb0[XN�@����(�V+fn��\�%ʠ���OU��NF��}�Π��K�!������Im��� �XA ]�oJ5��CA���X���j������&qws9����]7����I ȜP�Q5�5���(Ĥ�]
cl>���p58�>�>�A�hI{�F�/4��G�\�D�Ե��bA��6>k��!�8r�����m�9�YA`95=�Q���b��M8�MW��r��B�_��;�����\�m��OwH����@4[�sE����K�ڮ@�_�8_�$�d��ˠ�p*a!1�sf�F�Qڛ��-vA�XcZ��r|1/�@��	����o���!��6�a�C�y� ���nw�t�7�����c�}�0;6Mč@�Y���mq��҇?G�r���c�].p�^ՄL'`t����zc}�[zQ��5��QE��*������X�v�P#�%���:\g��c�3ed�z\
2���H�m���~aTL����M�"���l������nqm�n-�-n���ȸ�&��+YX�;��'��Հ_0=A��?�,�4zנ.(�Wa~���uN�g�BلW=��%�������6�u�40�X���TK�7��'�R�U�B�|��g������]g���~�����x�/�L�>ﲵ�]Ϊ�o|��h���y�w���.���GU[��6�E���Ӈr4���\\ ����_�Ԩ)Ȥ�{�	A�p[@�	�Xcs��V���e�E�on�^F��ïV(PF�g������%^a�F�3�0��9H�婸�&S�Y���S��"����G��T�$�$\}0�~B�����[/^�k�ޫpo9y$�{�W�e~6uk�fd�V3��LN��1�k45s���ԄIE=+T���'i�r7Ҥ��-�9���rI�r[tĪ��9�*l�mS�M>L����q����~��*�⑍��� ������J���'�u��	��131�]��|�.*�$cA��f������g�o�)�O�K3���bJp-��2�|,u����/o��k����nR��ۦ��7���)�Z:މ��P���A�Ǌ_�]BEܙj�p�
�Dьx�4wGD�˚�脱V�(�+�c�o���%�X|���zg��ݿ�R@/���a�
��,>0�?l�o��fM؝�|��{V|�yۙP=��&{\��R��:�ϧc�&����Y#�<]q�}�d�e���x�	 z`�����[����ϒ>#Bbt'�+[�[f���� ���a�'+)W��1`��/~�IB�O�?Ǡ;=|��?�Xy� �����C&�>�n�A���V�`�'^��}��lvN���Sx�A ��~�zn��Sz�r?�!	1x>}�쏠w_S�)����Rq)	}C�"��WZB����g$eoK��<����O�0	���7�Z$A��+`QϺjb���n�Rs�S��\�ݩVy[
���}�g�6Sh�'��J�W�:K��He�j7+���,���Oļ$��>�Ȱ�����[��ǽ�`B>m"����P8��W�υ,�ϧhbN}M(�� k��m��c�o�7ux�h
 "D-�FFLa@!�;r��^�J�Ryhh�∌W~��9�Z�("��i��'~[� �K?/]x��S�39����Z�(� h����6�h���4Ň������m��J�=^����5X�C	��
�@[[,�l��'���S�-�f}��� s�� Jf��	0�`Bp�o@L	妓�o����~�ڿ���9�����_�_�7o@��>K!ة�
��Fc�BQ���I����uO2Ri�8�wc�r|	k�#� U�߿	��'��y�����)�^�ӘBRH��	)��:���d�Gr�;�1�O�B->��;X�V�Ja[i��Y��u���]<z"xx�a�ғ @&�e�%`�q����d�dEj]�Z��G���3T$9�|mԐQ"�钰�E�2<,7�3w��O\*w�����p��'R?{�-Y�1��d!��N�Pk��TQ���|�����(����\��%z�cR�=\|wj�œ�Bxۉ��O�V����X۞$۔<��7��Fz���[�Q���DU���H��:VC���	L�ج�p��mJ�&�+Q�)&{PCS6Z��w��w��>?_���u\H{�2��陓!œ|9�C�P����S#7L�зn��nIsZ���';�b�?Z�-R{�j�_ GU=(ӓr[4V,�?�̦[9ۻq)�U����ƚ���x�y�%��h|�do��U�U�A$��>E�(�U1n�T�Ҩ�y��9I�`x�g�#T�0[�L������R|Ax��eh�Ov	?����(=����yU��Q�f>�(��t�v@_����P��Q���p�Γ��BjF&���zE8� :5�٢�JOڷ��ARb7N���~��1*Cj!�ddWq�U8��-�>o�-�8k(U���z��NgwK�=��oF�	�{e��"���Z-�"\�)3�w׆%�h���@�X�l� �C�;����$i<1U����5��:8� a��2�ʘ�}�E_�jtJ�zR���]d����F���g���''&E5U^u� L�iq�	��!���{D��������  ]�Q���G���W��A(a�_�6�>���A��F���J�=����oFFRά���w�Cn����3bbt�{�On����lh��>D�*l�p���~"�($�n��O�
0�{q[�	)O�)g�N���S�8n6�d�j�	vC��M�Q��8]�n�EA܉�R�㳞U\ȿW��`�Z��v^��yb�s0l���z�ny/;g*<@��~�$�_����P���<o��0��r-]�����EZ�� ��w��W>�*�
H�,����Z�ٔV`>��7�O�ӻ�Z��:� �x�Q�;���r��:��KxYD-�a-L�ys:�ɳU<0'�����ԇ}��"�����ֶ�����;��jߺ���q���sd@;�质�!��ETx���Y{(��:Q,��l�y����&�?�K��l��4�ȻM�zޔ"^�����~����V{OG�w��*���*���J\� ��v�ஷa�({�@�� i����������� kmf]t�W����*��#l�R�mC�rޏ������5�)J~�4���/�6*���]���r+d��q�U�x��gQ2��2a��l��5�X'��+�S%�K�(+���Pe�����d�zs�
:s�����W:�6��5�h�Dg����<#�+z�D�k�C�VJLHK��qj(��rh�gA�oĔ�����2^�x�4��&��EY�?Ί�<ft}�g7卓�+��}�xr������d�+�Sp��L��98��x2�Jf�٩dp�!�8���sR	M����/������E��p:SR�v�_�L���h&'���~��5��S]����P��,&*V��ҫne�Y���d2�?�z�2�����ep�Ɔ��`�m���.�x�|�����e/�I�f�K�)����=�~nf�ޠ4U���[��3�ՠ ��	�^f���GL
[���-Ͽ���1h�!�BőgP�F�qU�\�]ӥ_~?�#m�
�RT�Z���/Az=盡����ԣ,ǥBb�7�o�f�1��V*����I��L	h�Y0�N��_��⸓��)%;BP���p��X�`=�s!�
��i)J�N�����
-��3�����Ȥ+�k�7�~в�^,9���}u����5��y��I%����e@*�h^�n:����i������pئaq1�{^��
{ϗ�.	�����Ƥ��0g��� וX�:s?��w��;X%�l�����C�ɜ� Cmg����3G\]�S��#�i[t�A�Ϫ��Y��'��؄��" {,�yA��qqC�^��[�*�	k �	sX�w̸�o�w�h��޺�-�:��m7�� ��Z}�]��Ni|�h{��Jw0��p���y� �H�0�����m�g#3��R`���pu΢
ob�T�`D�Rw����*l��T���A��..x"&���b,���~�κ��9�>5��{;Ի�;|�8�'�YvN��.�i�^0��'x���������b�yFil�Hq�.U2Qjo&cPh�θ�g�d?W(r���g�3#}�ۤv[@�ķ�3| ���.�4L�*_����s60ɘ�c`��&��H��N��y-\����K��ݒ��y�<'�E���p�Uz=��mOdp'b�&�!�m�z��΅��r��3ң,qL�!�|+�J�or��5d��m!��~�/^ 'Uw� [�
ﶔ�e��k��_�<X]r~1�$,(~(<�2�DS�l"c]�TTM���(	<�yN,ti,��u!2cCTb��;̸T\S>��b���]�⚲���9̻�T-��{o�CgF_�1������Κ�|U��W�~R�γ���F'��g�T�)9X�f�j&���]g���rOv��XK������"�)�4�-=:ѷ¿G+K�w^��*�89����n�#@��o�Hv�@b�K���'�īt&���pt��@��iQ''�Cs�� �$��B>d��(��3��R_��䄗j���P�$�B�v�(B�U�5.0���\a� ���M	��MB~��)�R9#&o���.���G��4����J�=b��JYI��[�\T.�1�������¾�1̻U� Y.�NL1C�W��\�k�C�H]s���ؚ���D�x�ckk$F|l!8���yd�aӓ�eT��%X��F��j�f���oZ�N�AݸK�!�$��<B���އ��[���\u���)?m��/|_��\ �1�U���rx�s��g��#L��0լ!�7Qe��F�$f�#Z�O�Z=��gd�.��<��?��3��N���g�j(tt��i�&7��55X�����^�����H$��*D*rR|��mo[�[��q���O�Ĵ����Ήr����ZV%�ܑ�J�ʐ旧��JPeP�ĝ�'>��R�"��;�(#�H0D���a�!��֏�<1�9^�Z�N�߶B�8S
�<o :9��I40 �v�����W�8��+�
P�O��l�Um ��ϴ���@z-R�� Q6�� zJ��e� ��<C������?,�u>5��ٓb�7v����9��'!�1�Qk�'Ώ`>
v�ζ�\XCBI�T9<(1�ܑ+��F�*[nQ��h\�-�\a�����!�O۸�����ìu�2��6�>#�Y>q�/�O'�6�H����G����Ćh�	�����
��ɕ�J[3����(�KR�hX�*��,D,X�{?�k��) 䍍P�`+��ՠ�h�q����%�̋K��ч���Z��YN�e���U�\�m'��Ԯ�� w#���(�mL;���\�1��y�6���!�S�1vs?"y�=Xt"pL��Y^�F�|u�+I�:��@B��ym�.FZݧh'��d�i5O�PU�Y���og���n�zӕ�����٦�"����qnu�4M��)2��1ݬ�NI��$ �q7R���B��a�%�@�����H��iNeϭI�T����/9�5�7aj0��"�4�,I|?�~G���_#�0Z^�����V'�!�-��2�wDc��';�teO��a�nJl?���n�yјĴ���}��t1�c_�f��8<�}�\�m��jHۋ�Aі`��S�}��g��ֱ�����=��U+6�u?wiH�f��S�)g��!HfKG����Y��	��d� ��^2��Ԝ��� ���DD��k�����X"������3a�o��4ڒq����g�;#����P�T<3{�(�����b��od�m�k��@�����������5��6�˔>bO5�>9%wt��ൠm�$�<t|Қҙ�8
`b�����aA2_�I�.�n��k?x��{z!�����
X�N�x�Ŀ�������z�{���:�O�]k8�c&+�P|�3�5Q�e&$��ΆW�H����o�ǯ�����ޖ��a���~����O=�+?tZde`ʣ �Y�j�x[zj��$��H	ٛ�v		ǂ�v��kZ"�:w��� �Dm�B��lY�2�'��G���yg�r���Scq���*zp�/�qw��I��j���_:��B݄wy��ǁ_7�Z�Ǚ�6Oа��^e��{5�
�r�Jh� �o'J���~,石D�I6��F�[+�Q<��1�#�g:��?����ƜTc��y��b�͑�P�u����Y'\C��E�XVI�6�h��o˽DrM�U�XS��ƄiAW��f����@e2��PH�w��w�^M�=�ŗ���n�0����Va5�V�ΠZ������1W+� �YB����d��[�f�LH�{��/�@��"����.��?�Cu���{'�d��h8/�	z3���mPh%����g�=S1	�ˇ�`ѹwIu��;e\�O�ՠEQ��Y{��Y�M��K>��'�>�7�����f��+-�G���� =}��Z���kD馗��8�81��3��}m�Il�qOՅ�,���μ��v��17�~�W;+�a�KWe6�l3rǠ�5��O�6ԉ]XT,;�F�]ݬf�.K�;��*��lJ:�h�X�d�"HD˪�a"��(�i�SY��Y�Vդ͌�W+�\��S)[6>�,�mM��^�Α+��G�o��-A����9�<����1���G�3m��X�./��DM�{9(c�]Bq2#�s��U/��9�U�fU�ww�/,��Ղ�M�_���>�s�Yƽ����"��E��e� �*�_ؐ�r�,7�����3�S�+`0���#U���|v�>�H<bp��V��l]�xB���j��y7r9Ӡԝ�t��4:���9��tT##�<�kL|��.0W�^ly���	��Ş����+�Zۭ�;��ߵ�_�c�<���1�xa*Wp#�&f�=�7B�h�������]�:�!-9)�2�~�:��C�4ӒG��s���5��cq&�g��hm���Fd�8�V$�LC^�Fs��WԼ���ї'f��͜���y'W�Nz"�2��D�}��TN��pU��r�P:�`c�JW�}U��%�̧�"��8*G�=��� ����*�R#���J�C����^�vF.�o�J�S���5m��h�%��X��)�D�?��ǝ���L$¤������\:
2=˄�U|D	��E�i߃��Q�py;�yڽd��o�J�Dڷ.ߌ�����m����Ղ�e��:�v����\k�`��C$���]=~���Σ�ƆeE��#��"�P�����j�Ik��@�d/��99yP��J��B�+�ڽ�:w�c��]o0���g��U�c�?��ml�bاL��$�p�_��AF.!Q�p�*H�?��{3X��}��'��Ţ��i7s36I@�O�ߢg,~�B���ߊ����^�ƾB,�
�{J���&������������k��v�'����4_|��,�=�\���Ǫ��v��!0D8�p�Hr�E�p��{K�_8�����4tf��+R��_$2*��Y-�89��*�HRJ�k�d4���'��`��dj��zN��x��jS���Aьp����ߡN��+�M�e��cDtO@���F¼!@�-dX|�c��期Oky��d-vj�Z�B��Z݁F�P���^Q��& 3;
�H;u����#������e|�h����Y��
�K��(�}Jƒ'���J������h�0)"�D��X�7�XW�ԃ"��#G�N;m�t�M�`��8��)u4�!�#� mbb&;����!�t4�{e�g͙����,�;�j����5܁C$el�U1Z���@�=�ť>H�����ʲ: R�7t����r�X �u�f�N��Q,��D㗶��X�0Ny�9��Q�����Z*{=j�ل�&��%�0�P4���$��V�jh/C�9��t�Ͻ���eKM$���D&0 .�i ��MH�7�W�M�TA0|nu.M�K��d�syw����)�m����v����1�1�����9����p�zєA���Q�րu��\iP�:�]%R��X�Sr�2]L�{��F�"�ԇmƧc��F�K)j�������
z�L�L/N��y	:>ڇ^`���~��
h  ��]�9�*7J��~rq�����$��Y� �����bi����F3��;&&�����#۾̶�w���s�Pd�����d诶�%H철c�'m�����k�B�<Up��a�*eg�;
�7�5M�4U�>B嘌4v7rE�/�4���~����z�7ϒ
�$I>��}Ib�*��}�f6�ڄ`ԔV��[�)e��qr�yDD`:�w`ɮ\�I�pB�Ȩ�A"�1i��� �HF�h�?�G��2��λ�Mi(�9��:�80�Є=�й ���r6!e�}E�ǚ�C޳?4a!|��Rě���1���`Տ���#��O�?��&�Ӟ�MY�����	Փs��ktH �n���~E���9�N*�ee��Yh~0��K���M A���r���AY|i�hs�E*�B`O���º1ObXIr��8�/%���E����`��Ĕ#��ÿ���S {�Q>}�pRR�ze��T�r��G����M*QL��^���V�&�s
p�HO>,�RL�#q��k�^��fg�kk�{`�n�9�QB�?�]_���u��2�t�W�-[/�e_�U59[��8C�Ӹ�����(�/܀���R���eG�Z��n��ɗ�f�`r�̔Z������9-�?x,����l��H5���@Fp��0����V�y� Lc^�J�A��]�_���& �чX��sQ?�� &kg@
�W
+I$��2�ӶtS�%H@79��ˈ~<`�}�[��x��q�SLr���pn��c"�� t���.����}B�j��_�j��q�N����`��xǁ$�,����^s�I����M��eƏ� �Q�Oy��t����7����`�R������S�Rr]���Қ�z�����63C Ű�}��i4:�,C����y+��`��7�@���dl��b�� ]�К��$!�iJ�8�c"����,�͞��%�Y\�^ßb H�2�\��R7L��&��	��r�m��$�D�>�0��~��ڪ�ߎ���\��8�-S� ���L�3%�i���Nqn}9�}� �W������ߜ�z�OR�D �jt�HW�^���;��3�!�a�B`I���_�����s�b�UÁBQg�"}Y$ B,�t�#�I��B�=��K64n�O �L}uD:�_��#?�c��֮A8;5���4_�Ja���{,���A
d7�T�Jƥ}l��x�v���W�-D}�q9�fט�y�c+�K�6�֢�b�̚?�:�&D:fhAJ���	�Qu���z2��kDM.�:{U7V�l�C�s���������@�ڧ�U�;��e1����6_v���\���"xl��v_	r�Q���'�����~��&z_Y��.��.��:q%< ר����{Ѕ��mǮ��Wh o����G]�Bh���1��-c��O���R��д���H��i��N���S �"�T��Vz��Cl>=e3s�la�������_���&�b��_�y���H�K�j��+�D�V����oT�)0Ug͝��Q�=Cؠ��/ˠ�u�mQ����Ѓ��of�;Sq�	8 ˗yY�'�`�/7�B�cP�\���͎�oo{�'��[pP�i��}T�S0�8ˤ:;My�/�Ӻ ��rQ�+Q��Ј�e&a��!��2b����a��tr�ё��+O�����.�:*�ƖJ�ۋ��]W�z�u_&��E��4�p�7i[�y��iu�(Т� J�-y_i��m`��_)�j�_�Hd�7�RsV�B&/�1���țV��G >� X�^W�K���J>3t"4���7F�~�:$��U��#�*�@�
���+Ζ_8�-�&�I�f���,	�ھ����b��YՑ1x\I ���rc9/�$�Ω���2�Y��Rur�cd}F���X�O
%NZ�h\��X*�'����l�s�sY�z��G����ݤɰ�`�['Θ�)�Е�C�唌,�g�O���X�s5��
�ރ����!� �44�B�3W�J���8S6�c��Ծ�@%a�ߧ�J�~=(�]< ��n���ڒ��h1;����U�'P�=��1���S0B�'Wke��'*��:��F\[mS��U������� V�b,�A�,�K��#�])L������THb���m$jX�c�K�ʢ�����/��C{S�w?����;�k#v�Y:2ۻ��?$" �ۗ��.GNy�,u�cqQ疲Jt�ն�������Y��5<+1z8r8d�l�Չx6p^��M����xx��n����"u�Q��y����T�D?�g�9N&m�/=��C���8�<��?��ig�����֩YyZ�tI�HJ-��E�jR_�w h	��b�݈n9���pߠ�z/��~�t���|��k|���K
��gK=�B��� ��)�my�<�*��*�]0F�G���f~�;�̻�P7�E��K�g�N;7�5x��S�G��(�#7j��&��8i՝E�
��r����@�Ru'(;�O��x��r/��4B��#�lQ���KA���`�5��$�-N�%9H�v�Q�f^����M�!��a�>x,®��鴢�BΟ<�ңu!�G�O�H���F���8�d"������_��<>b��f��f0v���>�1	(�I��m/֢ 1�9�a�,����ʨ��� ���j�'Ԓ#$��MV�p����%;��	/��wnS�w9�R��HY6�+�vt�JS��1�n�kA 5�����κ{{舎�"?��t�o�ݽl����|���0�v١�W1�� ݿ���6M����թ��q�\�2��[;��oC�h<��Q[G}G�����
��7#p�������\(��K�ë�Br�PdF.RY<)�i�3u�1�&s�_)6p��/]Ը�Ȥ��3��:+y�L4a�֍�������j���::Y�����*�|����NG lR�$�ʑ0b��9�6�Xf�Z�Mf�.��E��t��8�������Dfr�K:ic5�aa���fa�g_�p`
{���2?A*�΍��U�q��n޵\����c��cB�i�Ajf��q�������d����Hҙ��������^ k�+��j�\��/��6��?��Y�3�sWzZB(3�pL�Q��U㑖�s/���6=�ż>®�ʘ������-ݟ�3�hQ6��4O)��
�f�]0�A��a��h��T#er�QZF�m<z������c?�ݽ}���]H#�>Q��}��S��{:��������+�w��lP�f�L�O2�)�t�ד�8r5ьd=(S��r&�>6�9&L)lB��\�^�9�7Vܒ*�v����7���"� ����d�����Q�*�Pq/
MF�52®'����w'y��Z��u���}g}	��!�Y�&Fu��Ⱦ���s��}��\��+M�>J���=F�dO��h"8 �n<3{&��X���|3�]ۈtĸ���X	�������T�����4om��r�/�=~9������O8�}�hߵ�8�F����o|�X�G�;¶�Լ�.��뺲r��XyA�H��4����<�\�;�S�1�Hh�01<q��Q��W�S�����Oʿ�S: S�wq��J%�klwz���gۡ=��p��hA�^�����U�B 8	zvh�WvĦ9)���=�8߮m�Z��-�:�p�j�������s�$\�k��>�"���Hq �����6=l0V�B�}��7M}^/;'UI��yj��/�9'(����cm���<���V)F��Yo'斘ο�G=%�rq*�-X�$�_J�a�<���>y�wқ������w-��i@� �]�z���4,�����>R��m(��yJ�I-:���nq��'w�8���2	��*����R���V�eg�C���}�U�&*C	e�g	/t���}ω��j��O��9=�,�,t���ri������f�"AV�^Ý[eK�k��t�ɧW���ٻ�C�z���KP�<��Wod/\�5����6qsp SZ��?F����}Wz���d�QH`=r�$�F�P=IGTJRx�[�历�^^�ho�[̂�CZz�+P��vWEu5�q�&]�͟��?�w���V] �����'N��l��m �9������.T�r;=W���5*M�U�Y�M���L�xM���ㄨ��PD"��7\���j�<N/�� ��Sc��`Ll;����%��B+�3'��Nt��12�&t� � H9�ʩ��Н��0v�msQ��fr�����C���h*<�m���Ϟ ���Z��@��66f��Q��4m*Oj4��BK/�P7~���8u�]��g��ŉ�rks�b+r�)Z,�|��σ�J��W��X�fH֮��@e���:T'���{����p��T�G3��r![��R{������%(�Q�����Y����2����}s�`�Q)`���@N~���ן�����꣰����� �G��N�� ��z?��ڊ�58'���a�>22
��4�����d���|�i=���G�5���@�pͬr������o��^���c����B�c���6�Kכ˂�<��������:�O�D!�K(#�y�⚋��M�{q����'?L23��z��F�b*�?fr�X#�}P�e�A���}&���7��nP0�Ď9���!�%1�bE���k�3�W����L���o�B�#s���@VL�NJ�xgQ�h��G4V~��K9��<V����Y�X*��C~��3��f��y�,*�=PD"ԛ@�T8+�
�5�>��Cdͳ��,"����ls�W��$���cQ��k��싶'Dchi��vO���0!�֕�EwHC�8����~�ل{�зyQ�պ�N]�(y�}�N�M���Z�>�ו�� ^�(Z�) Iı��._��B)6�q<Ǐ��쫨zt���3�r���Vx����L�N���+���î}ƇӢcZ',=ʊ���.�d<n�o]=��l�J��;B��rӕP�oB��|u�u�ƿZM�M�����՘Xc�(iz�6��c�Wc�xxf����6�&�Ԫjh� u�M���o�Y����}}&����|��[�[�]<owx֪FK�����0��-Y˵�W%ξ�f��QC򛎛̓.u2��V��<No��n�T�����(�����j	qj��@��hPm�`��~�
�B�#Q��44�8bsF�N��s�L|���6�c��ۨ�yr��>+�щk�]����U~������J�rapE�_��f����2�s�����<@�-g��D�SYc�'`c1��Z��aIU��l��w^��Y�k3u{���ß�ז���>�;V��WE�"�C�7B�X��r�Kr�P������]�(��$A`H���~�,(�U����n��A��* ��� :�a϶ͬ���$:��{�o2@���N�Gί61�5�ņ���<m�2L �g��E�����I	_�o|L�rM�|���
���Ǔ��e%T~y6Վ54�:|�	��u��9ք�z���2�Վ�%�R�cھ�ٔ�~D��}io'1��Y�w�Q .�Ť��u��*��!���7L�d�G�B���yPw�r4��?�iB0��4`�ǩ�
x�e����v=K'ex+f�	Ԓ���)�A��j�\+�8,�^���:9t�á����D5G���(�SQ[��:0`U�4�1��#�k�e�t����>�P9�	�%<�, ���1�y�v�������D�-B��V�R��$Բ� ��,$wFl��%���b�X�"l����:�Lh�nڵ���y�5p�<�qyp���b��y��GO�K���]b~c:�_9}�����Nb��%^���A3cnB>u�s��C/��k�H�{y�^n���/���؝Nژ;E��k�ug��J��Fκ������";�J��|����:)K�Z�G�r��e�L�ڙ�A�����=�H6"�ֆf{=��.q���Cև�%z���6�A�c1������u��#q?�u�e��"�Q���D*��P/�|ON\٣y�ސ~���T��u��c�E�A��%�;�JT�����?��v����F��ad��_T8�$��!���>������h�Ф�@k������GX�+�zw�5��P<ʄ����نmf^y�(Q��KS�'e�����\�\q| G�z�VT;SR��\f�qm.�&G)'�1q����_�1y��#N\�˦W��
�t\m4��8ZM�%6�g���-�~�yT]l��B���Z�S��2�2�)�����n�[��:�ʬ�4Kk�3�A)C�m��j��`%��]��?6]{����(Gi����نw,��%�Ƭi�+�5�JD��!�g��C#LĿܑ��)F��ͺS��Nt�V+(�e"�^��>���BvE��v?=a�NG�lF��qE7j�M.��!�h W���)��)�����M�o+�6�YΨ�����{0o;v�'�L%ɞ-�yNe
�)���FXfB���k{���d��^9z3>�k��6.z���'�n�5b:;��>�T��z�$�Ц�"���93�fa��F�E�M�U
��D{'�	�#�m/q���!9���)b���^��_�I2ʾ��&����]\��nLp�ۚ^c�y��5��p�٭=��.���"Z�b�H��U��*��c}�W��F���tj$�IN*٪G\~T8�#c!̎ժ�cyU)����Y�dC�z����0c88��	��Zw:�M
k�V��C��y��^�F�Wέ���E����z�=�Nf������)��$5�>��0�DCj�[�)h��e?�����Ch����Tn���c���i��8$��I��q�̀z��:7�}i��,`/�-����,e���A�t�(]\�@D�l7!�8)9��8�ڄe�o!{�.B��#��<*P�fl���̠^8�a��moA,��n	�W�7�Smh� ��R�p{�1��w�,	�yB	�B4^��Ŕ�6v@����eîh�0�~�?�~��x�`Fk�R�G2���_8�c�\��}����[��#`.�k�&��}ك@��฽m�Z}{�mi���I���܉�Ex�]���8�r��航&]��`���^���mF�{�ٕ
��G�D�tQ����ć�f�3�C���]�k:f��LaҘ{B�FۺGC ��E�1�7�8=ԟ��h)K�+H
��(���B_s�)��X1�Ȩ~�1f��Kt� ������̆�mGJ�1��T5����`\��R6���	�)�Z��u~�|� ��n��+�O0A�e��diZS�Ũ�.�{��"+��&
�F%|פ���Wjt����%gX���cC���p d�e\5/-�X�qz1��;�QIR�I���"t��#ѳ#����1`3�a�����Jq�P\�]��Q�u����A����㖗k�֛��]�Zv���ׂ�Y��ꨨ3W��#���2
��	]w*ȏ�Ϲ�}��S�>Ö ��ȃK��S/e���<�UY#�`f�`��s	 i���3���KQ䁉IBM{7�aNfXc>�?`���&�v�����VZ{�&��g?���,�t�ϵ,��uxÚ�V���[$���؇�S �l_��:�_���VF�IKH�IbL�Cr3�.RG�R�m��bOA������<�'y��q�p�_e�����쀻� ��*���_���
�K��usֹ���
�!o�ekS�h�2�������n�k�yt��th�������V��B�0@��[��3��=���mh��m>��_d��c��E6�� ���2�-?��&�EUt:�gGJ��Ru} 1�5Ȁ�3� 7�pA���_4����� ���K��f����
�M����q���n?6�����N,p٢˖�\J|�	��1� �¶�"n�E��>.�	уL�A5�w�`P���p��tb�(��]8j�����B�v�k�@ȫ�/@�_�����w�[*<�%P�hl�y�Tw3?*D'�WN'�W��"mע7����T�jp��\3�79���
�c��nn7 �*~r8�(����Ͷ&�V#�?����ݔA`{������-��r_��H3�9e����3H�g�]i���{�t�g�L�d���?+bm�<9���V��6@���|��]��8�F�0����b>!A�y�O����h��NA�`x!�Ģ�`l�1V_���A��z�~do����aL�H�Z�J��������jg�>5��� �����{��1�Q�5Pf�C�S{��&Q��w3��]�v��yVΤ����u�����n0mk�����.����eF��@�i"[5$�)��<�5��� XP��J;OuyQ�����juID7STr8`5yn��ϓ�˩��Ԫ{���!`'u�����0�����S+�m��#Ş�O�K�-��4�$)ɜ�[��ݥ����hǨ�gI� �iOC��MQ������q���)�jS��N���)(�ٿ΃gm"?EUzG����jw4���x�YՓ�.vk��q���[t�j�+'tR[��������/���z6����xf$a�Ht�*!Y�������!ܥ��Z�3�a�fzeW�+�2:R���\M<$�����ٲ��9:����7;��N�~����.q�J�`}�?�"�%/�ы��K6������%�l7�����DxT��u@	o�!�[������D%��(��+T�6�/9^G*���3��x���,c�}�%8�.=���1W�؏YQ��f�4�)�撁���=��PuZw�f�' >����n9���6�	��^�r{�n�]��1�pk�Wt+�k����k�q�Id��$%�*@�{d�Ay�R�Y���y�;�C�f+�0�������F�T��ź�Ex'.
z�H���Db��-B��Dy}��ۘU�FOq�$���2�532
��N$4'���U׾�E]x3���@���[=qwZdZ�~�K�� ��GcPG��M�w4=�?R$QEαNt���g�z?�Tߵ�5 "]��0�Ú]�w���dgб%u|�qdr	$:A��X<�"כ{��=�RbzIh[]ASc��~��'�5�{Xa��,*t�:`�DF	��-�k��g��R˟��{�a��2�^gA��fh�l���2�>/4�083D�*�Ajq�Dx�r^E��}h��[�j��B!�
�k� =ݺ�"��=uK�I�Y���@�sS�?�S T�Z�j�{�R�g�[��kk�9�\�_���z�f���V�v2�͑|F�5��P��	zr�<�U->1��gm����e,���L�gGg+�Y�y���'��nH�Jp�W� �-�r��HG��o\ �.7Y�����wn���I�f��.��|x�k�Q$�	�x,���$me�y5�ۿ�h�d^��3�Χp���$�!'�E=H�zC��*��=���� 4�T~���>qQ<E)��L*�eq4�N�b��*����أq�����Ĩ�ml����Q�H���0����"�D��鐋k]�*S�D�a��m��@I5�=ɥ?È�9��#a���ޑ�ܠ�o��u�I瑾��<נ�>9^�*m�8��9�*�k�]�ר��`����<)s�]٣IR�}��xc.
u�e����u����&�.-F��MHSM�;fp�S�VL���������Bz��jN��[�$M<0_6����ú�t T_]�Z����o�f�o�f���Gb7c@�G3'�У�G_rc����[�>�������Ԣƪ���V�)WŨ�z#��-�v�0e��],� z:V���b�M����4��&���{�����>��j���5����$�QJ����eۋ	�k�i� ����m�ų�Z����mI���<�k�K%�	H��8jT~�YQɦl-�:[)aN���Z�&�#s�d. zG@/w$�0j��Gì/�ʅ���\蘋T4+;�G�bQ�����c`n��z��5�vO��_AT�����u �Ҥ�a���=��>�a��;�,�D<O���J��'�c��#
]�#�K�� �UT0��D�Hy��?�}�m�4JZ݁��J���3۽ݲ�U3�y�w|�:����{@"v!
8������zsrWpo��Vߓp�rRnnnf�B����i�C�k441vH�	�bT� �g���6������ߜT�L�}q#t���;��XޅKO���
7����t����8eÒЁ�[�Z�Y�g�t�J	R��f�h��V�|?��*?�7�8��Bu�����sIH]�7T�´��O�ቭϤ@��w�S����3&������.�bu�s'j�� �Mh��61Z�VM��&T!�X/+�����aC��`,���2�읓��H0L��k�������1��Bp��ռ���	C3��b9_�b�9�ǑZ��'!�`Ie��/D-V��G��J2`.e9*�D�Yj`�ɘɬ����l�O2k.�y>2#�!�: u��+��hR{��|������V���d�T�t�Buj`h��0q��k04-�M����Y4ح�Ȏ�P<��~������8^Z �R�D�t
��wy�;:nm�~��ك�۽��@��T�$J��x�H�6e�X$�/� ���a�o���(���0�F[s�`������n�)�O<�J����/�^�yÇ�B7��5W���.T��岞���	��QI.z�)9�/}���ӇY�AMw�����U�# f !V>��(��Ocr� V?��d�`@�ܷV���>��*���~�S���,���h�h���4�OO��՞��(`��L�#^-��d�,q��)]�����r�h�W���3 $��p2i�Hb5�T�G��
��Oq��bߩ���E��7�]�(�$*��2��7��a��d����g���6ַs�w'�������J�_��(�O���T/o���_Ȗ�7�9��C�����f%&��~����60 ��i�����=3Q{>(��p�pF��3d� *��v��� >\��|"<r���e:Zt�т��s�������,^�᫣�n}X"׶�0��F��O��栮�w1������ 
���M�<�P���'��	�*�uS)�j�c5&�����C�%��<���!HU|L���zH��ܼ�Ŗ���0�#Z�? ���Jű����"`��s ��:�w��Kn��c͍H�2d���dK�<����`߂ډ�ࡍM�{Q�n���pF���*/���uC8��^b�t\+@'�u`�I��u靭��nJ>�)�V�����x���#L�[E��[�5@�A߼h�����>�ki��=��e@�l����_O��>&i��L6[@ɂ���-�~��x?m5@q8���I$���x_���цqOy�� e␚0bl$���/����-�)��'dfO2�R.x$P��j�>�\����;/��JC?ɕ\jvJ�������8��pL�ۛ[������1��Bn�̞�K��I2�1|�.78p�%�h�Îrz��U�fB�<���4��ᾊ���W��B}ȅ��~�:�N?]�s���u�vH���H+��UtM���#u`��p�vN�!��cJm{;�HԌ���� �F3�ΩKe�ϴ��#Nu��~�1��O�ٻP!G�&E�
�,��q/=M%rz�M�ݏ�%��kb �o��L�~�[�c�^�l�ה��Q4�b<i�^�Ot���1�|K��fp�a'٦(��8:�FKJA9����B�f�$l�t!Ex�7��� b�`�\<��}������Wt	��'��dWMG	h�=u8�O�B� ��pY��;�^��<�:)�:[�� L(5]���t���k��s�Hq�[.X�m
ߋMT�mX��yC11�x�	�M��I�wX�'Eg���72]OvX��H�i�E<jp]��f���Wz{WH<���ys��Zkb����p~+Z��͍5W����w��ϐB ����7�c��i+A6&�p/���a?��с{TΧ�����x�u�7Uǜ��.-� �j��i��H"s�J��s��Y����MJ�"��8vP�-�P�<C��$�?��ҽ��Ϳ'q�$;^�F�u�C���GtL�2(l��#O���J�|8�y���	�<1)����dל�	.W��d����(�c���uE�,\,޸���D���|��K��SB�3����;�"b!��5�z�p2��\�LʭB��|TN�g}����4ݸ; �Gi�6��M��T���p�Z_��'}A�� ��k��4g]8'��(U�a����e���nV�~\�|��G��$ f��t��:����[%�l$��t� )�L�pYb��D?����L*ʧk��5o�8)W�v*�/ p��1���K����y��"|H�JG�%��,!%��Ђ��_���;�9�!32>6�n�E�>"�����'�uݥd*��9�T�����fg>*/��+d� �ug�Jw��'7��1��R�d|__����Xp��.�9�a�������U�$�@�>[==K$�wѬ4K='�����)�M�H�呄b}�O<Q��%{�޳�"@���k�E%b�|�ōZ0P|�b���U;�iJ�'\�}*(��l�4m�`���`���s�\oQ��������D�5��lN{�������H�Õ,1�y�S��sF鯜3�-+9��@�gV�E�u˺Yǡ|��w�_z�u��l�s����V��.	�:Oq�&����P�+	0"�Y�ʧF_�m) -���n��SX�L�ֻޕGzn��5���j����٤'����G2_�^dT1���U���74�����j��݅D������`Ռ����w�w6�CZ�+���L��ߨ��(7�t8�e`̓e�dlC��Y��( P�	|�#��b`�5���j��)��pW�բ?|y�&+�0e�/2�Y��\�����җg�;5`���P|�����ވL��E~�N�]���F��Иd�X�$���ʶ����!����(�yw�v#<�y�Ӭ�7�d��듛�tm�k�6�"R�R��� Jn�ؗ�?���X�R�a��f�1GQ��
,Od6q.5�x���2F'�7)��5_EM��6'-�U�]R�:��	>#���ɔ_]#�,�����Ó��+�`׵ޙ�ɦ�tj+'�aR�t�c��f3)3��hI��pY�q-�_X=�:��1,��p���;�	E������*%��B0��]��au�̘��{��wݦ�T���JQ���i#����ɘ�B2�HZ�iD8g����U�G.���P�Z�y�i�Su	�{�*RKi�ʁ��	�,� �
X!M�C0��(���nO�!9�o�Nn�lq�$��Q-orB�N"+ە��P�C&-s�C?�U�H�����s�I7�<�N5+�ʪI�c�Nk�\I,����Z�=/�C�s�R*OE!_-�&���ٵ����dn�L��g�7&��U74G�ř����v>�H�6/5+���~�p3�*��1l����@��B�1`�e�0�!��LD��]:��Z����"ud���<'�`FZ��MD����iz�C��b�x��׈�{���3-Ǵ�A=��rh��Zq�X�}� �m#�jo�?DM�P��*�s4`�Ku��r����j7M�N�@}m-���U9ؾ1��1�ΰ�8���⯞���M�yp��1n֒����=�����p�p�*hF��`f�?��o^�J��=���[9�X�]1Q��r���'� N3Y��x�j�~%�9����!1d%��i�X�:��t����O#��5�n8*�a�@?�8j�B��q�[ ���$�x�ٺ�p��L�D|b[ �3��hJ_�%R-/����CN��Q���.Ob�^�EU���ی ,�<sܳ}�y������X<h�{K$��&)�H[��~�I�c/)��A{�la�i(��b�ҹ�9է��Ӧ�^�31i$2Wx*w?�|�!�`�z�E��&_~ܫx�����|Y~�Q��uO��*��_�2a���M�_u� UK��Nŕ|I�6�X�Z���o���wrװjڇצ��
7Y1�����kי<�-zع�<>�+,�m��[�l�zZN����1d�a���o�2������ݹ�5��ul9��CU�o���O8��9�]z� ^W?]׈�x��am��(����82 ��G����+�H�6��/�p�O�Wp5 ^��j�x���պ�B��FH�Ʉ�g���d*��ȸD�Vs鑲�f
/�"I��Pt</�)�������랴�a#��Ĉ�RmׂUs�0��ш� "4+viZVp_zLba�Z�a�
*G��a���*�}t��5��[�d���}c���K��{#�p鰺q1��_��eD�M?�	Zv&<G&��&c�7dK�X�6ď����_О;ٿm�\<��������A�`�d������}���*�s���1�������#P/��m��T��n̛(����ϊɴvZo�K���,�s�6x<�&����4J�@ԇ�8S�/W ��Kr�qT(��R���f�J�}3m����yB�%7��SaY�K��R�1�7.�b��F�3�X����1�͌n��^�5 �J"EIub�<tx�[���Q�2��`�?���1Y�x��?���ў;��Wjj.�ץ|M\]�Y�$|�!W ��AއfI��O�cb-o3���yaR�{�9����w;��}
+5��s?�Ϸ5-Ip9 !<L��ɩÒ��T]6��JOmGh���p�����h~3NÅ�?���=�l|D�/��Ra+��2��ļ�PC|3'�����#����s�ey���.�"n���6}����߫;f�p(Ьt6��s�t'�2Od�C��n�~Fl�y�uW`TG."g�@�q���P!d�ZXM�S������ �t�n������Oΰ`��*�n��B���Y�?q6�bӈ���=��c���D��̦M�ښ1��M�\�:���n��
:��,�>�Lh�j;,�I]YN�:t�5�s�(Y ���rjl�8 �O�S�Ć ��L���
 �XJ����M�ț+�1�Y^�n���md�mG�g ��i}ZP�7�����2_�?���,�w�53g� �)� ka/U��F�|n� zL���?Dt۸4Kgȃ�u[�77��8��0�7�LֈE$�,��	UBy�
Z��2񥛅E��INCP|��F!�Z���l�f����f�l��������q�L�u�#G��w���_����ך�aB��Hx�5��S�tɬ��3��������oyog�a�]�0��Ԕ��&^$-R)`� 2�Ϯ�0XL���\:���>u"�ķa0d���s�\N�R�C�WLV��<�/X�ļn�G��~,���_�&�K�!Q�+�z�,��)n��p����ު!C�
�LI�Λ&�F���0=�u8�7@}� r�+6��YPZ��@(�`� �ml�d|0�y:�U�Vh]\_��=yXJ"���DŠJ
"�ԁlSW�M�bѨ7cz^�S
�#1EX�$�Qi�����P;���%<=ӓ*�ڢ���	���5�ܨ�C��)?�o�!&w����M��1��m�䟝+o#Ƞ�1#+jb�=Y�͙F�����R`1���Nb�{����J<�k>���Eos���B�q��xV|D^����M	"���w�y��j&�ͧ��5���١�$�Q�F�
J�΄�=<�p��`���6�b�����K*+̄U|ԬF�Ӛߚ�����
�^>����\��?#P�F����rZ����U� Yf �rr�1O�����jL�\�+�$H�n�-LD��4�i� x��M�Е�@N�vL�e/��P2@�a�{
L�ˌW a_�;\�uIk�:z{V�t�B&^�xcE���@��3���n���KR�Њ�D�\~7�I���C-0o-�=ѿ� �!������]}� Ig�&̓�V�6e_���"J-���T���0�U��v6bq�$NZ�r���>��Ui�bu1�����&tA���C@�K��^���H5~X��|yo������ ?��к���ݢ\�|R`N��D#��l�**�э0�l=]���ڬFGq�+I�����Z z�-uEA�MǴ��&�pߚS��M�Q-��
ϝ	�o3#2�O�������7�;��Y6�;��,$\혊�c���}��u�'�����VXn~�H���]r��4z>�Y<�<��`�U"Xjv�i}���"RJI��k�����NgNZN�&��7O �!�DA�V�7u�6LQl�9�b͗��(qKCW�����e����n��L��5���XB��I4-o�s8-z {0��ؑ.e��,��S�,�E����ځ.�k�5��*MH� 
B
��E�2�b�Q�%�����!�c����I	��$�u�
�W��J�¶VK'
W�Z〖2��㣋5?۷�����.���X$ć�G�Tx!r�ŗ�a#�+��%AU~zݡ��.
��R9��b#*F|VFɰ�i�#���/;sY�4%�4e9hŦ��.�8e�]� ����S� aL?��\8��Vp���]61��ĕ�8�>�R�(�Uَۨ�؀$��&@u�40J�ԧ�_��Ϛ��-Ԩ�f��!��u��'���f���XS9�)s�v+��h<�[p�����Uӳ��ΧD�3��Bq��y �c~��B6����9��`0��rmPPp�v��� �,�[�eHႌ&������f�0V�_�(ޖ��m����g�EqMǕ`��Uw@�!{OE�3f?|��z?�j�� ��6�Po�����6e�s2�*+n�k
�GPj�[|y����n��F2�2U+�0��{{ڀ y�co�q�?w����,�#L��F�����2��@�O"O`�%-AĦ��T�-�K�j������簫�+��HRz�¬~�z¹�As��a�q�#�W�o�0�tΞ69\_N��!|L�c�m�����e鴤���j��|.���/p����hc��|w��ik�< |��ޜ��8Fw�1�jN�͑Z^ks��]kT��̓j�A�@6H���.[����~�a⤁����d�-��^���9���&hr%���b �Wu�'�l˔[�b�a�f~T����Ri��LB���-Ĺz�����A� ��Y7�?�02��b+���R?f%s�5Kө�(N�\�)����G���gt>���DrH�N���2��w�����s~K
]��T�)e�X��w>�8�K�Oe����&�L�+IW��~��(��w{栌���BP�u�c�O�A̓-�*A�4!l:4µC<��z,T,��7zi���X�G��"��N��
-)��(����9�.����[YW�x��E�_��=�BU��*�sG�״N�&�'��1���\�	K���=�i=B��G�%еT��r������Yrڼ�#i{��0YW2
GjIw�_�0.��n<m�c�5����@�$cS[<��<r��*aͤ� �*����G�v:�j)���+g���9kx�k��r���N-e�=�؁jܾiiԿ����Bw� �k��w=��.����Zb	�-�}��Jx��?��h�
x�r���zFlxn�p	��*<g ��e���='志���Y�>�ճ���'�#^���Ǐ�q�������o�,E�	d%���Y�a��@�~U�DL��`
wӼ�X�+.}Z���`}{�_~�+JU���J����s�h���rL���Eԅ���yM&E���m];�a�JY�������ee�˱��g����v�iY4>A�Rs�a\夝paa��J
!+Ʋ���
�`Z�f�A�lʟ��t��[�L+론d��ĸ�zD�8p��	�s��?$�-�Y1��Y#֖���ـ2�hq��)C�q��MF��_�X��UZ}-�1���9[2����E�ҁ���:fj�5�(���*��
� Il�I��0� �Hdf���[�y[2�;�2�B 1��ś�zE�ƥD���l*_���`�����_��)5-�N�Y�d
k���2@��w5�j�F���w���8ۉ���t=T�a�>VdW��F%(��0��?�O?}D��?,MbL����W����$~����ɒ27�,T$	@,�)������r��hm�����ɗ�=�'
s0�gpNיִp�Eq�ϣ*�
6D�x���7+�Lލ"5��$@R���K�2X�eQ��0"�V�G�������7���B{����l(PĞ�C��|^;S#�Ȗ^D�l6��E��KJ��~z��f�L���IW��f �s��7\�jEB���*ۦ9%�P���A���sX��O+��V�Uq��A�
(��G� ��D�ǚ����?��/�お1���"�+!��P��m	�WI�ղvDg?��Mu� �)��a���6��V��^��8���0�����Ύ�䬻:cU����6L�lw,�9����jz9X5�qo�E�����!�&�n�7Kp�&��|����]!��d�2��V�n�=p����,3���Uh����oӃZ�7m�
r�%�h�s�v�#�z(�1vxs�iص<n��s���}>1}�#9'�G0건��p�� �\Hw���T���d ��!�����v�=��S,A�H?s:E��N۶鏶3�Q2V`�v�a��|��ُ�@�'m��G�Y\��ތ+$�eQ�ؘc���"�r��{.KXc`?�&��
���6�|�hn4�_��gW��?�I|�K�S�V��c;-n%r �.U��M�e>�$?���il�L��>]�A�tۜ��*hF.{â��1K��њ^2x�������>��4��nT;�Ƙ���S�HWͼ�X��%�(MlZen�Z��˫ ��&�(����΅}�V��!u]���HAvl�K~]�V�y%������,М���D�<��J���Cй.���B�"�� �G�aR�dt�R|fz	���^N[a_�A�V�H'��\c�>���x���4��[�PoV\Y�X�/@��c&��p��i����A�?!�Iذ�'va�ቬ�Ժ��y&a�JR�8�V_�r�5P���he:��̌�F�Bm[�SǕ��|v��t��]��w����q�(F>���7����֎�p���U�]�l��z����|u=S��]v1{����6�[�B��(���Zh���M�XBl�$�8�f�v)^�x�����+�{�⏓�8��/ԗ�j�8j�C��*A8`��=KNwM@8���z� 4������
Wu�<����V
p�չ�oqϳ��Sb)oT�Ŷ�j��-�]0��q�Zb���[:z���w<�����H
�[��0L��Ϻ��VJ�s�=�r��7�J�~#�Q�	�l�X0��P�J�`� �ǔ��[��l��{a�O�m��9�;���0`��p,�\����T���p*���r�0�|�,�M�I�BSĖI���J���h���9�v��v�� ���#)�����k��s$�q"Х��oH��]񊇜�E�ۮ��T'=9-?M�]5x�*j�'�����s����߫Túh�N��ΫF�&	8W�v�kGde��'2��7��K���@�v韴������z��@�C4�]ѵ��(�Q��CB�sWE�fr���#I�6]�#(fݭ��7ܔ�yV���'�  �i��]w^�̵�����U�d0����� ���+��@�W����0�*M��x�g�t�Q�\#��3�C$�-��8 �b�I� j�z*�C����ȭ�C���3�}����t֜לI,:%�t��0�d.eB�zldi����F�nWG��Xmz���v���$�R ϣ[G7��Ƚ��H%��;��y��w��T!�W��;z�B�J`�xA����F�0�M,я���e�m9L�n;Na:����<M�Xx����farS�볔���84�+$ ��:����m�Q�e�M�s�HU;OB#y�l4�*ߤG��	��l�n�8nH�g��8I?�-�M�½' 
�q� ����/+'YÛ8p��>�զ۔�E�~U�E����3ݳZvh��H��ު~9���0rc[^���|��9��l�N�cfs����ƞX77Cѻ��6��Q.��M�G��/;I���7�o1�<{�.=ȝY�	ݸf{K�^^t��.b�U�5�3�K,����?�_�eJ#�4�N>��L�_L�N\[����*E�bH��* �%�J�A9'�}��)I����!O-{�f#�,d�W��%'/,�.�1��7{Cx��pD�n%�M;]�ǿ̫�M�1��FV�C��b�f�q��W�x�Zm�S��]�s5�B�����d�r�ۂ�mP:�����*˛tL[�Pk�/h��l�S$��R�� ĝ�Na����H��
�T|�� 9�F���������MѥQ��0�y
K���d�a�c;xf��V=]h��0�?!���2HKQ�S�gb't>��y�Mzt4��R5���6;�C~�W�2^�Kq���~�M���(J݇�9��;c�Vx���,s���YӘ:�kx��AV��U�]��ɨY	��о��B]�eF��<���5�+w�as���Ҁ��9��!ɿ<���h��8y�=�B���S����'7�Yj���!U<L�6���Ȫ��Cm��Q1��>�zO~>|\�j����:5Wq�ٞ���H�ۙ1K3H@״��[�fU����ހ��� |_:Q�OL��z��1��M%���C�Sgax9���)?�0 y�K~�>�䢯��bD�W��&�1���i
jZ��������FG�r�Z�]��ymz�[͘�i3p
���l�*z)zy�Q�~�]ݵ�1�ZMD^����� +FK&��h�H�A�&o���p3V���&ιm��/�K�����-�g����0�W���?��U� ��7��I)Td���u�m�*UK���9�!}�M���#m�;4v� �	�%����В�hg&�q���}Ċ_	w̹���CI�B_,�D]��%�m5 �\����U�%f���� D��g����d�u�#x��?���Û*��~lJ�(I���Y)?�$�V�8.̱3�[�&��10�sp���(�L"Y����x��URj�D!���e�N}v�S��:�:�mn��YEq��Y Uｼ��ߙ�Ufk4��ƒ�-R��^�cb��B【��A�B3��":�ok�P\*
ߔ�Ҧ�~j��XhU�i�Ǥ%\����_��
,sJm�,�����:�ʕ��[yC�9U=��`̺�M��m�$���֕ܐ�[1�ɑ!�.z�Hj������B^_�ggpa�u�+8l�r�'LIӗt�C�'ɺ$����7�~��]�����a���:<���J�{�R��
^=|�J��h�
A`�c;����:�ȅH����˘�)E��p�6��m^�]*�i�@ �O/Ћ@�2�dbl�Yѝ%.����W�����2�#��Fb]}�"����[g�,oX��-������yzJ i�!��^(�g1P<BI�:G��m�`��"o:0���,��k'��Zǡ����:�2=h��wg���l�Q�G���[ZA<�}|8/��0Yx@�q�}����a*�������u�4��� 0���\��Q\$��t�ƨ�P~
�,/ܰιY���;]$ucQ$�Zly��|��
����\~G��G�JV�4J�����K|�W(��w�r��7�v[�َl���Z.�Z �/a�a���.4�F����cC�Q+�W:�`В3n�x�u�-�R�=B�ݛ�������5vL�^��?�I�d����1��;�
������ S��89��р
��<��|Q/7������ ��x#�?s���ǶU�N�Tg-=�<ٝ7Q^�:�փ��z7)$�� f�*P�u��M�B��zfEj��Y#O���Uㅖ=ЙiW��}D3���/c��̌�8��<N�򭼥�X�ׅ+��_g�³��}�2�y�7�E��/r�Q���s�T��Y:�,��6����-�L�J:��/��$_KB#1.c>��I�	˄�6�N"���zuL�pے�Us��}`������ջ�u��c��9m��92�ȮQ*�>b8ld��gП0�Ϙ�2mA�
�ߘt�%V�e8��}�Pw�`ɡ�͠�f�)��MNo�i�����~�n�%`iܠ���1�� �����'��:�? 7Rc#� 9�ma���E���=0H����L���~����H��N��FEv	����Ϡ�>U<	� ���c��v��J�},@Ҏr7��!_eɷiW�\� �lk8}�5��Ѫ3��F"7����%-�!>��7����K0�M��K��?�~�7{ac<�/ǔ��� ��`�0;�|2R����	?��v|�+]:[N�$��B�0��1S�'.O2�@�%�6�|@g��i��(���8��zK߱�M�D:7bD��������q�㚯p�{�?l\���H�%����6ȁ�h�����p�	v� �0�x3���f'�Ma�9��v�����۸[�IRr��pun�7��G n� v��m�����O4�i�VCk�F6p�.�2�0�������E]�!E*KefoR����!���u2u�݂P���&/��z��N�D.�U.#�A�Ύ9\#��*��]�  u�@�Dձ��G���ނ�׉a.Z<�_܌xz58D������̺)�k^ �{���.ck�u������N��6�9�l�jA��� Fn/�1��M�yz@�N��5�Ǎ�ЏM}\x��9z/��+��Ge�e(؀�z ��&wX�?��E�A#}��9#�>��=��멊��U�jI�SA�7\�?g��J��C=�y�2���ma)�x��v�Y�I+�J�D
z��ti�e�����@���f�q��C�1������.Z�ѯ�5ίC�(�����_!�����Vg^!�5�v��f��a��NO��C�h��E�� ��E�@:���!�5�N$���I	R\7a[g��RY��_r�j�αt�8�Veq�~0���]k\�s�F��0��L�z�p;��g�3��;�#V���tf6��
	��r��mN�(q��� �����a����8�o{e��7�8�?�go!nY��w��Z��*V��YՆ��կ_P2�-_ߔG���ҩ&
"L���[���غ4B���`R���="�NY�g(Ե֦�pZAd(Դ�����v���2[�ma+��r�F�پK���Ao��-.*��8�io�X4����dJ�ί����Q%|a�Δ����q�9�d��	u�NЭ��9js(}��)��<I����B���2G��*���@����\��{
�@\��D�,��RB$ P
�Uva�v�_L�b��O%~S�uf��Yd4�7���{���L���#4�z�Y�W� ����Βg�\�	`&ݛkq�?��m�i�)r��U��)#P�M��J���4�;� t-IE��o,�=U��&̢���a9���5�B��xJu�ɹ���-[0.��K"r�R1=�9��WH�7�r�fȶ��%�"��1��lQ%^=�{3�O��XZ+�qE���<Vb�:��oRֳ� ?�R��"w�/�x�jR؝�匯��i�^"dPnkU�Y}�H��g1�sY�}�inx��xJ��Z@��M��X.X�|�f�ts�-�����o��;�tS�c':r�ʩ������j����%I!��r�B�{�3����SBjٱ�v2�m-z�7/~ w1��@�o(\۲��E��e�p�>r%ʖxK7��'��	u���y���)7��s�x��FA�1�`����K6�y�0��̱�j��2E�4�y2�Q�ZՐ��������Xj�f��?�]$������ܒP�f�*e�jbo^|���+ʛ�N���ji��d��
,Cc�N�i-Hh|���z���E�˄��Q�ۚC��$�e¢�U�+�C��޻J�*C� �8�=��>�>~����y�y�l�J�oP=��.��&v�x�R��O��|�82�8�{s�㣀*�傏m�>�.��2��]��l�kgW��b�z�nS�9�t��g��aś�v���d�7mCAUF���3�.ÿ�P��]��,g�O�`;��)�O����N0�H6�^"�ǳ�U4��"���8Y�"p0��;���7�u��ŕ�%�7Q���ܘ�}w�z �S}#�I��#�[�3�-�f����҆�Ia��ap^�G��@Y�����~����U���ҵ�,��VW���i@|������YԳn�ծ�"����G-��yN<�WU���ڵ:�d.�9� �ba��7�d������9J��C�6F��fOfA�v�KZ�<��}��wԛm�,��n}�����S��I��;'Y$ v9�fK�O��S��AF�A_�~�`r��32>�'����vof��347��D4뺬����,Jm`�1�~+ד!��")6��Qw ky��%ؕq���Z�GmM_�7(��fQ �_��@�ey�Izy�+W�W2U	h�g�i}3�9u���ϐč��O�r�U�޶ O�o^OjREO##��t?FRa�z��O�7VF�{��5\R���XC����Ak��j{����6�u��s�hn�{x����-8y�-8�h���!�'RP'EV���u���p9:����fT��	���N~��c�"�J�M')h�Ri������8�+�?�4T��lZ^)�3&����V����8"��i< ��Y���Xx�}_{��hk�)��R�F��"����4�7,�ğ~���ZU�x^sX�:ť�~��(iA�4QԦ��N.q!���}�AJu.Ȏ�
�)��
������`O�`P�eq�s���m�܊@�=Ǘ�|�����S9�$��!�1�QW����8�
�����������G�l�F3���-��1�g���J1	��V�8��<XЇ�*��Ƭ^����vJ0/�3:4`A\Ca�<�K���6�\���T�|4c�#V�z8���姐u��P�-��B��$)���c��
 ���-F����� �-sb�i��O}t�6)p<�?c���i�C�	x��bӺ���ۺzH��D]H2@�k���V}7-5�!�

�l�����Kd���рa˻�ڐ�L�e�O�Ȫ��g��>>#� ����G���9qD��r�;�p|H�zj�30�KL�M�J(T������e>U�wK��.I� �����>���?�P�G����ҙ�QH�v��*�2n,wb��ܬfoZ�D�b���Y���֪�q��6-�P���y�u�2��4�\y�]����b�e��jD�\�0�q��� �v*�lS�N�ș0�p��ۮ����B��:TW�:��
aB��X�MS��3p����e�Y��5�/�%���#���ؐK�������WB[���� T	}��h^�m���VU��sq���B��9��R�ڼ��$H��o�x�|;�~%��*�OU!^��6������zl�����
a+.)�$:�N���|�qҵ���"2�
qQ�+Md%�0Re<i���ܝ���6_��&ir��`���|��?��%�+� K�?����(��5ܓݸ�U̙aVu2[����+F��ښ/�5��r��2�-�d��~7�L�7�ۦ���z -I����v�[%z��~�O�x&�s��!�+����f?(n9�����>Ղ��?YP+��@*Ϳ�����ާ��J�c�h�JrWP5%!d0dˮ��E��)"bܠ�c���9���@p��N�w�%���3!��.J@	E�����Qy
�t#���=�UIX/]�Y� ����͐]c�������v��j�d��+ �����92$g~�!F՛��[��Xy�����P���fF���������|טh`, 0L�xs�o9�	qi�����蹼��zp�������
M���+q���V�5�R����dmhj{�
7���G,L��o�S���r2_~�0؞͔R4]�^e?�O�a��ߍ��?!��5��mZ|��r�x�k	$\E�{����n�&��E��"tN� g^-��{�Cw�4>XJR0c�z��C!o�=\�]b�Y��/���y_9#�tCWc�JL_G�P���d�~:����X�� Q0w�B�cD�q�Y�X��qm�̬����v��	���v�:�_n�
��$wr�!)$��>���S���b�O�̼!_�UE{���%�P0{�6��ƺ�+��>T�h_�9	��g�.F�vn�rF�i8����h1;�k�q��0��-t�o���=� J�`�d0Xw����1����֍]���k�|[,���� f�ޠ��I�U��1�4��n��;G���/���MFAJ�J�α5h/;���B_���}[g��a*��aU.�{����/�!s�Z���@M0����F��Abk�ۮ�V���R/����&q�Ϡ�(�ŦV�>��R#8W׾�.��ȸ|��)��}݁Do���[;(��f�|���x�����P�G-� o�ٽ��^cQ�4�U+|,v�(:|��8��28>E���CRO��U٦c�%�s�5�A4�Ȼg���:��Gx��wph����w����4��QV�rC���������Dz%�b�Q�� ^���Y�`��5��t��>u} +�D?�y'N�_���tpK�R�{�4����Cb3O�i��:��ͻ����q��38&���`��U/d+X�h��:G�w0f+9�h�=�Ǔ�K�'֖P򐪼`tx9%������H����e�<.��ϖ0�x�^�u}ۛ*C���5��_�:,5H�qX���CPYbS�#J��Õ�m@b]�yM5����2t0 �n�����7�"}\�v��&���ǨM���aP$=x�1����j�w,{;L���ܰl޻=���GB����l�T�j��̽��N������S9�
�����Yk�һ��B�(Z�?z�B�vbhl'nr����\=�
�YY����gv��W��3A�?gΠ���hj��:��	 �. �s3�dS��ߋ��/HG9� ��%u�+t3v`Ȁv���xL�CA2®3��+�\B�#v�V�3P�'ce���
sn?]L�n��C�f�T�e]y��r��}��;�O3c������7��d�s���I��a-�rOF��0�X�W��`���"I�9MT�eS!�����z(��Z�ho�.�t�悰ڕ�8�_<��j3Ι�=���� �-�gm�[$�%�]"7�=+� A�_Zq����8X.��|<u��y7܌y��X� ��u��u��<��`����6r4X�M�x�^�#u�Q 6�+��r6����:�0��)��{AXq��7<<�;0$`�T��|�^��w�%O�3u��ޞ�#.��[s)dB�E���r�I���߻.0��lx��O_�J�/���	��z�k<�p$:�CLO�]q�Պ�e[�)�
�j������1�^��V�H���F\dr赊��O�����a�r��d�ടI ��*���8���S�;�zG�u�Y��pL�mD�}�2eK�l�M>��[ħ�LP	���������Y\��!1~�˥'��٥ ���Rzzv̙�~����h�45Ěx��q��vuo˫��?��ݮ�G�y��?S924t4A+H����뾏Ibx7L{l2�r��n?�!� ��*�z�JMD1��&� pTP��� ����zN+�}g���o���ϐն��lX�
�-��<�'�Ps$�vo���+�]u�7�o���\,Ǧ�6���{L=��4����gz-������Y��*�"��X�/DBw��-�c��`Ѓv��n좊'�#ßj$���`fQ����BME�,q���`BPOϡ��	�F@�/5�hs)���w��(Q�?Wp�m�Fb�Ag7`����y�ҏ[��-�2�e�޲�e:\9.�L�\�t��xo�A�"���n�{hk��E��1l;����}LI�_����f%κ7��h�Y8Q⫅iDuf�LIzH3���&����fӱr�?a.I��0$��r�Ub-A�,�Ln���������{��D�>KwC��L�li�
I�Iq��bŠ A�'�_���?a�m�D�Up��/��2��I�1��uo�e���w�)�i�봙��:�٢�w�ؠ�1C�t��0���?EJ��.HN�}����6��{�a��@�&�3Y�^�l��%�I�Kt7{-��Hے��X���:s�}d�b��P@?L����q�0:z\9RL�\��<Иµ��r�����[��K��>��
�K����T���`䓃|�m>("Z�ߩ��s��'�O����YT|w.�x:.��nI�p}�I�y%%.��?^e�=�m�{
�Vhy�(�m��[��u��y�[Fa�VZzڿBX9���	 O��"�6 �GD^B�P{E�o%�ұJry�;�RX#��W}�O�������sx!�uΌ�)�V)F��阰�ᴗ��"j�1y��jc��p;7�[�i���:]|�.��s�/�2krT��U�?�ߋ�U�w�	0b��l��wޑ5hii���Ў�K��/�!�9hi[a��m�+��1�� ��wTf~*'���ɓ�ɢ�8˫���j+�cs���-f��_�φu�_���i� ��!��Q��|� �}@����r���wsͷ0�X�A���J�����Y)���n�~�Է A|6r�
� �0��ojfqM�9��Q����m���'{�j�b�?�.˺X_(U�t�����)]�I�^ܦ��'�����gJ��K�K�oq����*���-���ZBva4��ST�u�C!-,ZRѶׂ��^����iJ'��;�_��pS��F��1�*��KI�o6�k��y�ɜ�%�3wuΈ�
hI�`*o�#ӯ��7�k��	�(�W�����:������!�6->>�j����g��qDh;���������|�us��ŭ"sWV��A���@���£�U�#}�TQ���I��Wn��2}�́��ۍNG�����f����o����v^�d�t���v�Rj�u�\�Q%)G�����Nک�
�y����h�C6�U�@��Um'�����a[ n��;V���Cm['�9kP���J�T�:���Ex�}��dW�u�q�d��������X�FM?���vI�>��8�_���7|�k�`�۠��@HE�ܓ?�H^/e�͠|��鷺a`m���p{[�"3t�M��Q��A�>�u�g�Aq�E���vQ���z��Z��N4Vu��D2�'�rZ2�����G�Z'��]�K�uɄ �/�t/��_=�g(T���ص��۔~�fK��m���
�k��|*����z��@����0^��H�{���N�Td>�j`�PD n�L����83(��Lr �n.�,��2�65�S�(�ś?,&�H��g5(���!���je��7�S�2�F݀�����z*��o��+��?갤�k�,{ ġ��{OX�%Rݝ�R�[�#���A��5�5���&'t�=-��Gk���{�Q-��U��z�,�x�`�P�w~���9W�"im�#7P��q���.�y���uDE�x߸����6)}� � ��#����t����/y��=eT�o�
'��*�gᩰ�{���61��{&�W�|3�!�|�����б8������5	����C|`�8�)��*N>�1M�m�����ۼ��~�a�A���q3�"" �:,�On�G8r7�V>	�Rԭ��_�m�'l�w5��|~�Ew��~f�@*�#��	5�����ĺ��Z�1�r�Z�	UMF>� �J�^��7'Y=4��B������8+RFG�0�����Aȵ�+nV���T�2�|Z*��>o��5���t�A��m�[�Չ�����R7$�]�y�ӑ��X�� I��='��)�_ �n�π~�<���2h?�9�t�zx�-.�Q͠W+RԘ:��~�L,Zq��R�B����̧�[K<}C�/��Hf�X�QWM�aRB@��o���Մ@���ʷ��J�pj��+|���n��(ݙ� -��g��|��D	<���ILƉc0�3��l�gZ��.Q�Aux�� ���+��!]v���^���fc�4��n$��)�v�PC�)�Z�&���V+~����uʬ��n$p��oS����#��<���)0�ҡ����j�5Cq�����F��Qܯ���d�Z\Q��Z��cy��R���9p��i���-�S/�k��`��-]=��Ŭ�oP�r">��m$���M�$�ScE�V�ɭ�,�Yj@������y�?'�m�w�E��?+�+DEoqd?8����P����q-�"n'�����W���j|lr⧴?$� � [Y2�67��7yZ���j�=���	���a�<���"ޓa�e��'d�������ΰ�{ș�뿣�����pDN���I�ǰf?Ec=�(₇�&h�9M �t,�ࢀ8X����[�f������2XB T����-%�v��dId��ah=z����K�����o�3m��ԥz����m+m�؜4K	��r_ϫ^;y��8�N���:>�kq��DJ�$ۢE��(bH]cFl(a�$��ClyIJ��������u߰؆|7�4�	ڭ��f&c�ߌ �M7^���>�w</Դf�7/%G��|�Wp�5����A�Dr�`�mx�S�Y|.��H�Z��k�\�/��&Ï��Y (>/v���F}�fr!��F���{��D����p{���K�O?�g�,�o���-_�ٳ�x+<im�,>�V*���BQ�'�Ӎ,���ȍo�̼���Կ��[E��/�\�����pA��U�{�V`F1٩�n���8;-��+�x�پ���A�����Ư���6m�d<u}S��/??�?�����(f\(�U�2%6����4�cGj<DA��1;��i<�e8߰ ÊE��n��vb����&"���L�F�cڴ��@w�2'�� L�%���1(��g����4����/'ZU���TC�<��w`��y�,L��j�)���q
]�Ѝշ���R8;�D���`\��*�Y�G�۳r�J�969T+����w���[���8O���fK��H��~+ڛ3�������s�Гk/6:�f/Ҫ)�p�L~7��d���G9��)-3��3>5n9~�2JP
�Љ1h-|��t��QQ%�]�.@� �o$m�t��ш]�[����{��y(���2e���-w��V�y&}�T���X~����0uF)p��cɧd#X:R��qV�p���
�k�),�Z���9������L7�c�=J���ޑ��V�����(���^�7�4�yC |z���K�����?�1]��Q��."�|g+�:S7�8|0�U����оQ�M+��X[�w��˗ ��_���(3cM[d]H�69��F��{�!��w 3������&=Ό�0^�=EU)� �U����\�4�0^b�u�<�U���-�5�O���iB���^|T�_��pC����u��̑+�nM�*�S',�����{�=9��J"�Bc�=@v��w~]�C��`C����yƿ�T��ԏ���gxI�%�+��W��m_UY9�-\' �D�dt�h�@�xl��h:k?ZK�)�~��������E��3�Xʓ!U������c�AfQ'�&�	��/ׇ�^�/�^���Z�����ñ<��H�\�3j*tt���q��2�����,�qט�Gm5����cI����1���ذn34�:�\<_^c�#���9bD��C��DzH9&'��2�L(�ZBХ#9:�8_�!i)G��,G��93���F3��5/�t���SL��u1c7�4�f�2�|Y�`��sn��oup]9_2�^p����5떀��y��6��Y*Ŏ��gt|Z�S�{W$�Ws��k�q�a��.�#�K�\h_�Z5-��X���3�F�'�`Y�1px<�/pvd{���Qz�Z���6��s��)�Ɗ��(:)�y0�#�ɾ�U�V��n�_�f��u �2��sr�,sK�K[ zΛ�_NHF�IR������5X�u��+��g����$�����*oL����'Y�P��9X�"�e$ز�u�)P쒈~�W<͸ ��Q��-p�%X]�	�!@4����X�"�t��Q^Ls6��v��ry}�Rвzōٳ�~7��BS�t��%��n~���L�bY�5�FZ�c �P����r�����!�%8���9�X�sI@H$c�b�Ȫ��X��*���דϛ���q�m!lGrtud�?�a$-+o�.�Y���uc�贇X�8�a�QI)hf��[5lNi�{����p"�f�S[qD ���s�����FS��[���������ںnj�H�d�B�\����8W	�������~�g�~��r���]?���~�����Y�܈�KX\޺&�*��;װ���%ɹ�G���m��e6L!!���M�E~F�+��Y�KՌ�a�`]$)�Z옅 �(U��$�g<"�����PV��̿K$� �cX�Ǩ��8R&��[��.י>8��2��z4�"$W����Y,��4!(��E5z�����j?uG��c
��ȋ�d+c�2�!����(͔���w7tv=��Ύ�Ԓ�ݬ��S�D��W�S�
��Kdpz�0<�ڏ���l�����mx�U���&�Ss��ө�X,vk��<hab��mxk�}�e6$��j������xw��uɤnˍ�wCi�bD���+i�!�۱3�a�����`��!Oί�y
�
�[�!K2�1���Gۯ�����G;��2\�����bH��1��iȑ�4�]ԕRR�����w���IЂngG����'a�o��W��n�N+��5h,:�ِ��ֈ��&����^+O���1��U�-*��2������Z��ƥV76.X��,��Ǉ.���kX���/���xa��G���7��ǰE�ی�wl����lu�9�xL�?~XG�,���ryiS��mZ���	b�[�d�!�9���8�8�����jj���;d�e7n�BX"�l�����D���鉖$IA.V�3H��!t;��/>@՗9�s��.�m(��'�sD:q �\���.IKyw?�7��cp��6����fG3��#D�@>o��T����8?��_�մ�X���(��Ց���Ȭ	����4~̋J��UE��bq�2�����oj5$i�Ŧ���3��r�tM�64~x�o���Z��LO�0aP�3k^�d�.���Y��Go��c���H*��wg�BS���!H�4-��dߘ��y��u$v~sɤ:�i�@u�J�$\��"�?�iq��\����%��4j��:όwY4[I��U��A���h? �$$V6Ӑ�I��b{bIW�D�ê�p�9��.�:J
L��#b1�.��˶A,9Y��
�VW
���/����4E�p�.+���߹�8�6e�>�R�9�X�O��� �������}������g*������jg<�4�7������P:TNƆk������oZr���RF!U��$=-��]F
}l�\�w\���g*��Pxͪ��^@���u~[[�KV0���@�S�4���z�w{/	��.:�Jؗ& �������]q�!��} ���w�'���$	�m��&	@�dw�Tܯ.�hT�Huɕ��6��
��F`KP��)/�"�h�22h
�B�h9vr�f@·Q �������YG�'�n0tAˌ�g�3�,��u٘�J^���eս�G(d:{�ɝՁ;A��vS+i����JC����}���TM6$r!�y��ba��)���Lu��o�yd�Ht�f)���HL��1�-��B�aJ�iL��U|�D3t��;��7����M��|{Z��0�n
y� ���Ѥ�M����)~�������!L1�NHE9��E�Gڕ��D����Snb��@! S�ޒ�*��*"[�G��w=�����<�%��u��*�W#fd!�M=�!�	����+?̠sYh�N�� 3[��]��
����	Z�ב���}�L�Yl`ZҗD�>@�3˺$�r���*�\�E΋ �%*擦�ҧ5d�P�ʌ�Ο�{�?�,�Po8����~����Mq���"ulAKR`�2�:��ic �D��8��o���������?=����8H�N�t���<��
���7�9�.�v���i2�: �)��h���V�W�`Bp���~5��S��Q+U�O)�O�a�ۡ�۽$�{g��􃚅���Z�n˶�b��d��J|i@#�\��DLf_~�G�[G� E�p@ψ���'��V��}u=@����^^
�;ц��V�+۟"q�OQ	�lZ2E8oM,;*c�9*i�z��:į{�0)�q�Ã�.�<G�0*G��8�/��1q�J�E8��tڢ>��Ԉ�/�M�D��Qj�Y��1��k������Y.Z��gѢ���-��*u���ڜu���vnͣ����k�*��6�l���0�_aѽcjU䌾S�5��Y�c����t}w�� ���5�o�ڀ���]��bw#�
,$��������pՉ��jwu���oO�ua�z�d�%hÆa���V�t��y�(l@K��S��O��)0@ďơ���[��ySv���q;��-!&A)V�B���1�d`ǆ_�c�sFMN��űIJ5�߼ZN�2�����s�l�1�;W*��sT��(ki���b�XB��r0���XI�+�?p�v��9o]sJ6 čј`YK"��#'��\�x�
���/���v�Sb)t!����?+�T���r�i!�%,��u��)��YSݷpK-aŪx�}��8q��Eq*;��Jp�x4gR�[��pn5g���u���������Eh��{:m�:���<Q��^�䝷>,,�ڷ�zxwFs�d_�/6!�%�K_	��m�0�U�2lB���&W��n`��T����T��yAF�T����h�:�nB�8�7@O���qmX�.���z���a44^m�����a�f�E��`��u�x���)Nκ� ��g��F���K9��c���%��Ƿ
���ѯ"8sw�����|������?�lz����&�s�����*G1����Un�m,>~� ��]�2	��Bg8�-���Wܬ̇�o޳I���-�KX4��������4f4��!�� Cn�Z�*<:�u
��=�H�N���������h�|H��x��=�K�I<�_�9b�$��y;�����<���i�&��^�_��;��<�����8]V��Z:�9"��6gF�bɥ��V�ގ�{�ѯ��6/�}�Y�v�؈e%[8d;��c�yYP�����O1!��q����7u��.q2^�j��D-��8��}���ZF��+1[����Kv��.��.@	�DT(����M��/k����L���}ey �Å���@�m@����(�)��Jr�>��x;y2�A02�,!��9"�*�v.ڴ��#�v3���4�^�<=nbgh��O>�K�a�&�x ��\�)]g�=>�����>!O��5�dˇw��$�r8Y{|>F��I5�[*p���<$8�0�5���Hk���qk�6�̘�&��+b�����7�",�hZgo:W�)̷�E���"�S<��0�w����Gu�Y����4��	1$�}�<«���܊�*�~@�-@>ba?��M��b��`;yL!������2����޽@�����~Ye����ܳ��;�RՖ�`υ�$���&ę�S����Cp��9� TLV�D:S�jP�3�m_71�<PVD4	�&��=���\|���PPԸ�����ݠ�-��Y, :3�&��`��o�mh,� [5$u�-�OҬ�Ek�2��>HK2¤Xд���h�weE�`����S��H��"K(���)eg����%�>���"DU�`ε%-�3Ј{n�r ��ˀm��O7�	�S��h��TL�ĈWNvg���{
Me]��@�(I<��yk���ٯƼ�I�?{bƙtO�N��/�E{WE�լ~��1M�Y�lLE�$�R���`�ǿ�N��)3�]�<��G�oȜ9�)�Q��?k'E��uƋS̤���%�햍9 L�������z[i�=�������E���C+�Q}�\CE>t���8����C��("��:7?�0�l7_DX#VG��(q�4A+�6����Fb�%�s���+�������dq·y)�I'����|��_�u�	V���+NɎP��7"}O�e�(ԑx,*�ة ���?����B�	㗳�Uc�sH@�ʇ�T�%[e4y��CևtVC�4����VprO��ۛ�/�= �(p!�����f"�Upa��A�h�nq.ō6�����]�F&p��44ND��q��Y��o�������(7�^QTH������B��uiF�����QU�$׽�#8_~���XāZd���T͏H���
��Q�BO�X��S\�т]
���g��]�
�vr��X��lp��X�+���(���z�-�M/�LJb���9I{���ZZՊ��V��d}�D߈�
�� z(��Or� ���l�T��FK��`i	I}����\[���0[KUN>EHK|A�&�v^?u��ɣ�3\ڥ9����	��q�����?M(�
}-�b��?cR�(�ף�m個̠��E;�T�x0��a��������[�*�0,��w�L�Q�SNKK:X��4���GB;����\�o-��-�#Ӎ6������NSaYn�M��9�'�����c*R��/���nW\F�ɹ%r��W��i|N�R�g�	J�X���g�\�J̇��b8�$}oNh���f%ʻ� c�t��2]�)FSq���2��A#��)��K��e�b�����M�c��'|[�)�e9���J':��ū7K�2l\Jf�K3�b��n�tZHE����V��Q��������1��V���I���9�<�Z��.����-�Qz�r_�v�5t���]�T?��J�K��2�Qf�k-4؎Ĩ~�ju��e1Χ������
�� Z���$r]���W^�^=��$�~��[w�I���Ti\�9m@m,,�������lP�#XN(4-߫�����%�b'�[��٨�%r���Z�����+���@�3�)Y���'�in��eL"�
d-�T;MGӐh�{�y'z�LÊ]��.��S�w��Q���\��7h� (�}T�p<:f�[	�}<=��z��VD�3v��2E�.��9�q�C�RlW��v�����JGwݯŕ�Q8v�S� �����?P���ma���sh)L���Vju?ở�v���Mm�~l)�����%)>����z�V���X�^�!
>�>a�։��(���<���
M%��V���f4���Hl�����ʚ>P|r�IO�ha�\+��nE��Ȑ�Ё'�ds�r�M}T�F�C�}��K�8�8�ٮ�x:wi�ׯeȨ#4�U!o�}�é���h_�_^1��)�ϩ�e������:��eՆen�0�� |Iȿ$���z�.;�Ì�(�`���0b�� jV��O�N��@�j�nG]FA}��M:<�(����×S,�!������]Nc'��E=����xN��v�#� ����7�̘���(�
�?�g`��fK�=�6��:���S�N%P^��J��݂�R�Z	�q�>�K�7(BF5E�����䞍_sˑ��5�b-+�D�I���1�����3��:#�ݯ2Ws�b2�=#g��WlՌ�Snj���I�u6���}	�u9P�W���~�(�.�rokZ E9+'�iŵ>oym���*��R�6� ]��Tz��Lj3�,jwál�+}����,V�ȗh�}¥D}AL蔢F-��Ĺ/����,�F��I��I@��öL���bw���Zj���0`�J^۳ޮ/�������|�CB�0 \y��p�p�j�Ƨ��^-~eײ$#�b|�Skt8�A����8e�y�MX�$Q@l7���rn�V�������հ4�c
A0�tMP-^	2"ce��/�yӂVX��A
 o�px$�
K��q�A3{�;��㍴;n-��<h��ئ7{��&ɒ;>�PP�KG�܁~^�g��`NZ�Fե���,JRb�h��ӝ_�0���f�{���[�X�/�a����rJ�����G�]C���춶/�0�h�,s�Y�_}\��ʝJlO�Q�6P���D)QPXv9��) �;��2�]U��\STzU��g����[o���1ya�0qo	�U��e���<���zc�ۼ�A��,(ʚ.����n��F��Hf�a�^%���և�����H9����ZO���3�.�4�ėu��'�]r���'K�sYE$Hn�+��� �����]��'����5UuR:I
���j|�S:R��<u���fø�.��8�\�Z��ړb���ΰ��XpE��:��Q�a����I�кK�]E������7�H*�]�ΏOL����)�γ�gEiP�_�2	�/C�VA8��y��n)�W ��>�^~fT��#^�i��'J�5��۾Bpg����7znl9It�'	�>g� ���s^��f��~d����A�u� I����=���pp�	מ !p��8���|��R���*v{.+,�(E,I{@��:W���h/��RDj����8#�]�U�l�Ԗ
C�)gђq���A���'z<W���[X�S��Iÿ/�����[E`���~<��o������1Ǝ�a��-x��$V%���	D>ɜ[���E����?=���_������lI%P<)5+���%��r��1RzIq�6�m�%���k6�n
8oW�CА[+��0��Ca�\C
h�g�pk. �`�X ��54�)�Ļ��J#�q��$�D4�]Bpuk'�05֤��e�~\�%f�ςT�PT+���ĝrlIh�Z/�/�o?v�(W*��צ�pN���H����e]�*��wҌ���7�:�Ϩ��c1����S�m���8hb��Q2��K�(�c{l����L� ���Y�P�UEU�+�����L~���ȿs���(6���=
6@D�>1!p7�%�,F\��g",~s/�.�v4�qD���g@j�0M�B��lF9�8�"f�5�2����Z����5��+F�ٗHb���D���Ae)��T�Y�~S�S�D�Ě!V��a�F\�m�Oc:���u��q�V�Юw�.��;������`�o�8>k�(-����3qj���3	��9��ѝݢi��,m8��
�ٽ�j|׮�%���l�*ID����x�l3MA�:�W�!��gY��.���lf�P�ShRh�@�~涎��B��D�,'�DP&k�/n�۷D6�s�MI���\#PX[�'��M9�� O6T�N�{��������Y)I�)G����	%�D�)���bВ�$y*��S��9�������j�����T#z KcZ;�m�d?������  �Y�"����hk �.��7'qǊ�E��u���3^�@=U"�$�횏ޥ9v���*������7�pJC����ХS��5vQ�ڿ~E1Mڅ�xSǶ�v�q��=gN	��L��#����?[�Ȣ�ސlc���Q�#��
�4�Tb�[ھ�����{�[*�B8��u�C����9fsw�����_��B����^�#Ƌ��x�0�闗\M��I�b
��~,��E�kcŀa�ǕJ4RW{$ u� ZU6��q���,��a�1E[Po)���}�C�r�q�9��DI��������_dZI�`X�f��+Q,�ɏ��%�L�98�`\�֏ܨ��oe`��/���>�|-8T�N�L���D��e�0�j`�|5�Y���@���˃����f��4�
�4c�� �o�[x
c:�@m����z����t��G�&�b� db�:���ʞd$\�v���.ig���Q[�7�|�x�qԿ6��U����	>�%�&�	E��X�s��h��&��Bl�cO�Kך��{ f-a|�%H~#` �1\�[��Y��y�a{����=����
u.^�!os�Z����|�c�+�I�q�{S��ڠ�{,�O�A*�w%Q9�#���D�n����ia�2tW��VY�����_���ٜ����0>��e��!Ku�?0��QO�C=RVx~R��R<'��o,!yL���~�����効=�t�S����L����7C56sg��/f�E,\:�y/��<ڐ�K�?�WٮMJ��ۉfc@e>J5Ȫ'(5�
�k2���٣�7�\��z�}W��c�@&U+q
���lΊ0�����~��Ұ�~����/��xb��|��@k;ˤ z��ir���˴C��QE����Z�W�7�8���%f�M}�>g4��h��vH�VR�w�nw��-F \m���+xocv��a^�3�f�8+�1O����9/MB�N�A�7�W���x�7c�f�.��3���`Q�^�EK�I��\���n�0߶`QIuZ}��e�Q0zVR}�h�A~��� �z��"���I���~�X���J�S�s���ZH|n�T��/~{��R3c�@7&�3g-�(ؘ�W~�a�Y9`h���@0%�β��R��.�Ϸ�	XCJ[��r��[�/�@3ֱW�>�����t���v��:�E��GZY*/J��P�a�����P�.	ޡ>�)0�O���AP~�m=�i��eB	�$hM����6W=Է�3�T0���t��{9�@�pN�A�4���@k�f��n��Lx��-73H�s ���ʬ���|��1�0�[4�)3n��w�*=~ �u۱��d��=]ɋ"�	V�����������s��߼����Z��	�4_�v`�J�1��l�X=6����FF��{����Iyz�����exXŇ�!�>�9o{��ȑ�<���/|z��(�{ތ.����H��o�\yAh�A[j����pL������اq��t�D�����//�Mf	/T�/��=�K�\q��13�uw��}ߔs/V���*6B=�hz����k6ʏ�r���y� �����Me�P�S{}��i�?⿞����Ӯ�HXO�	�����c^zf��<)$���2%����}n�Lz>~*�w��z�H���"�I���Pc�xUT^�۞9��6��3�y���;Ik�\�E2?�Zs@5����8#��D��a��.�*9�`Q�����K��>�m�X�,,\��uj��/b1L��;����� K�1P��Qi��JhK,�n��?�#���,Y�>��EGps����\}l���ʯ�8�˛z��`L.G�.� P7��e�
DY	��"W��j��Kg�� � >�S�L���<Lx�����X�帆�my�S����#g*3wv^�nQ$�j�7&�,R[��Z���q��=Aҵ^���>�2��1�%�ӱq`���'����*��nɟв�o(r؇c�V��G�n�����Ix��/��6n�3 H��u*�ާ�����V�%3��46�Ҥ5gn1[V��
!�L &��䆛������T�g~:���o"���n��_�M��]+�=��_�2������wW���7�#������ �1�l��H?�����"�UƱ�Ot���p�]̓����m4bI��UZؾ��.�~�9c6&?�ۉ?��2�I>�(��A�L ֟,e����h�z
�,y�Y����{�4v�5M�?�����ο"[�%�a�(;G� yd����ˏj/S�\ܘ!Lӊ=0�k`.(�?��~� �ν�YXt����0���@���Q��dN��v�����CT��`%���r���8O'Ayt�͟�X���5F��A��  l�0:]�����;G���[:���L����)��bu}`�>��5 ��~����	��[�즙�gec�v�T]��/�ޚ��V���|��9zDLF˺g�GJ������.?N�r���@��!�?w��0��;����N(��`��}�X�oݦbR�xi���e��i|_p�t���kys�O�h���"S��Q�������۸ջ�'V3��԰�M�	q�'AsqW� �<�h��k/"H�}u�^,L����*����S.+�"��M��'��:A�O��9����Cpgc��� Wݮ
�|R[�N�p��Tt ,�=��8�4ߖ��FtfVr���	��,Y�@<k~�<��]H!�eJ�P��e%��������!�^1��X���$G�����*C%��ť��f�,d����@jߘ"�X(�8N��j(3��v�ߝ��p���h�p�(�@��v ��W�N��� �L|���e���#���< .q&U$dP��P;ګ
;b���q�0B(���i1R�V��S���;Pp�YgـUA��e���4l�`�����I��@6�8��v�-�@��5�]�/�s]��O��+ G���{@j 4C���I6N[����/�uTK��"Q�N�P�r��˳�SBf�������|է/rt{�C�[�QQi�9��y��:7��q ���
E�Q�v���X`Y�p��F3J�c��H�Jлg��d���u\K���<�J/wX�r@_%`���W���Ft���~���*��y�+�y���2�g��g|{�m��Pe�s���А��$�݉�%]U�T��!r����\�j��v�� ��%���*x���x���:�����SI�@� ۄ�C����b����J��E�Uiv��ڰy����o�
O�-5[:�6�}�5m:�ׅ�MJ����0ы��p3!��(R��T2��,2�6C.k��՛��S��"f�	;�ʢ`+�wsWK�S
egRJU~	[.p�t�j+�8qB��"q8�`�V	�w�v�c43X��	�Q�֪�i1�m�r�#{m3ob�&4�.�H���S\x�5�u��|�i���6㪅�\�H� #qi��䳧N8��G}߃�Ya�6��ܮ��P�2h/z��Xc��UĘӌj����W}I�t�a�Z1X�mǹn�p�-�g�d+`8�����-�Rf��`��x�JM\V�����a�4�6���-A�i���e�z��d* �~
-�T��̆nMy�Wf�[,�)r~��=$�zN�N��zVz 6���bke��#ω��H\
�'��i5yn�u�{m���Bzy�X��bK?F���1���]֘�Mk}B}>):��D�j7C)�GY��Q�#sd��+������T2��˕k3OX�ᢙqM75�L�����@�/j�3�	���P7��e?�`�+)=[R����r4����i��R�V�����(������²^�@����.�R?!CHP9&�נּ�:���!�>���-M�o@シ��b����}�������-a�w��ĥwT���}�:�W	i�f2��yH"Q�j�*�3wc����T�n���+�&�S0d"�d_w|*�kq�D"���4�3��U�ٵ1�t��& �r�A�.���|L��c>N������,��y��h2#w�e�P�ؓk�{k�8�q�t�Z΄�k'�GJ"�VL��.ᶱV���}�[0;Adw��"���P\o��Mſ��]���##e�ƍ�1�	L7 X�V �D��J)�@��jO�¿~�����q\!ts�9��C�y�����u��)r�,Hlt4���E�SwIm�c�ڕ��JB�˷���Y�4cջ��a�A~�!v&k�r���D�����9�(2�r|���h������y+����F�Q��ԿM�x�v�f��ݥxOZ4>-��9�Y����ʘ�ގE�}(�8"V�y�%&��L�il�7����|��*�*)gp��L�c����8�/��sd��vՑ�7�g���Ulk�'�F/l� 
��]����)#k�T��V���w����?շ&�W�9�E��0��Vm�՚ڲ�&'+��TD��@Hg�C�%`�`��!�&���<֖Yy�#���^q��GS���I����2'B�G��zi�,:��߆�F�F�yC�z)t%��׉C�f��%A"��-�8��k�Ē�ߊ�[[7�1��?E�����H����K�v!A�O�L��бz#2?.�<N����_ĴK���X����F�d����u��"0��` !��>IW`l�i8�r�l��@&�3^��	&�0�4i?���42 '��)h1I�K�����f�a��ۥ�`��1�L�WGv��_�a
���wc��=��}�U�ki *�*���b���*Mƪiި�F1�3IgW
n�Jm���'`T0i�l��)�된����FqlM��=e/k����7?�^9hi��ˡ��;���w��>��5W�!*ɘ�c�";x�:���j�1�#�܅8F���l��lB��y
�qN�C�� ��bǜ>��`At5��-V-�4��g�L�����!������g�A`��| Q=���s���W�+��ְq�D�������'��s���N!����<�ܾ����p�Ǽ�/��c
��o��Yh/��W����e��.�4wF��Q)� ���7��D��n�&캬7p(���`�Bهy�]���{�_t��s�&}UB-�
�a��j����V��-=�]g�{���y�*��-`k>��`�{��%Hk��5�����A5�3R�<j��)�)<������Yf��Dz�aQ����z�tLt��c��Z$����Hٺ�8L��
(��k�,��OW'��}��j�h��n�Pޤ�o���*�n^,i8�	sǇ�S��6�)�I;��؁($��������5��9���vb�Ր��*�3$�����g���dt��xHJ�;��]7|1��F0�1��|eՏ�Yi�+93Jҹu ���E��������[w~�0
j�z��"��I&�FOw�w��!�*�BO�E�kQH����y*"Nq��k}\��cj�E|\5�l��
{��/��t�I����Z����e,���Ɲ3��sP���[���bU�P�0�g<[8�Pw���;=JmЊ�"Qp~��[;��[���N���4�� 30�N2d��d�Q�����(XU�-@�8�/}��cT�T|��j���h���Θ�$�CFmr��Ś>�i�/���9-[]��@to�6�����1� ����}�w�  �;��#N��#��wZ�"���FT�^k����-ia@���L-؛�����i�(jn>>Q��ED���}|�2�y�@)��{�_b��jG�_�}�.�̳���i�5��C7�̛��c�O2��4�.��T��������EUj�"x�9wM@��C���c���~+���g�!(+�������I�~$9j�ShK� �s�!&h��!W�L�<�g�w�0v�;|压�mu����7�LJ+�I(�`ӶGxpYiUC~��\�Z)��u:U�^ciJ)���IS 5XZ����i�Ѽ�њ��������~��)6�d��J�qB}��k�>+��y�˚�<a��&�7�!8�dd�H�,H'�~��(kw�.ḭ�/����B\?*�6�F���0�%�M����,K,�Q�M�k���׭,��	��m��pw8;�p��z��9U��vx�vg4H*@��^'	h��=��*�=[G�)�(L���r5���&�#�1���/��C!�HԵ��C���1$�Lo�Af�_V�c�ƕmE��\�Y�Kɀf��Y�w/�t�;���7YY 8�Cx����j�i;ؕK)��N��
�_����q� r��糼d�;�vA�{��1����Uq���һ�����m=bF�+��,}F�&�������Sz҉�lI+�ù��k%67z2��o7	�Q/�����,F�K�j��"�w��HV2�]�"�/����Jdo�N���Ðc�7���υX�یư�7����Wh.&E-+����[��n�^ŉ�f�u�$�1����Wf̊���kS����G����5۱t��]�`�,��$��tp����-;�{�֗oF�45d��Ơ�veyq�9��Oٳv��N��~$�I/t�K�U/��U�h�cg`���[������pʆ"y���@�*�Ad͗(=	 �I!5�F-a4s(~p��^�7�+Gc�y.˱�x�ZE��U�Z�����:� ��"�e�u�p���\[-���ż�΍��f/�����fl�V �f���V��������6n��T(�%w�5� �$5׍
��q��Ա�A�up4lE���Ve+ ��]ZJ]J6u՜�+�	m�jg,�#؄4@�Z&�;T��|��h̜�zk���>�T>�|e�Y.�?tԸa�q�Ɔ��m��<`�Є';S���ӊ�St�׮W����s@��q�c��b[�c���� ;���h���0��_Fu?I���A̳�<����j5G&�7�#Aa�'���7��w�@�t��!At�R�_��[3���c�V�|d����l�2嵸���j�<?m���3��C��qڐh��G�[�Fwb_N��[KU�Xs�����v*�,������%�6�;����m��˕M�k�_��%��q�k|���4h�agu�!�!�f��3��ߘ���Д@��1֣U�ߺ@[�VF�������H�|]��f]c��U�^E(���V����K-�&���e^�&j@+�J��  ����-O��?��Z=�rz�GRfoC<�������+J�I��Y4�	:���dT�i�$��� R_��T�I��AC�p}7�����ito��9^D�`�hԕ
�m,��k^����M��N��tC�80rsg��Y�wE~F��mцA$�
�{�3�% �)�`pgY��71�*L�YP
�_̍�w^b씧��}�����u�,�y�O7��4��x�q×��uV�����x&E��r�ȵ#���&u�HAaѷ�)SS�<��k��j�=��>���c��� ���A]�P�$S���u�R^�l@q�Cd�<�?��33i��!�Q��'1T�cq!�y#&�%Y>�	��͌*����ÞV1W{ ܈���w�W�r��Ƕ�͠vb��IUT��V�S�*�x$}�rD�"��~�V���md���W1rF9���x��n_D�0y�Y���9JZ����.#ٝ#S��b��5i��(e!�w��'&t*T�KT^�D��]������},��7�M��;w�1b�~�yG=�����o(I3����~kJ���2;��V�u��=@������{ ~a�* �'���
��j���r{/(�̱�E�,*�2C0�FvR\�'9�p�1A�G��Q�B�cMڐ������,B��/}�d�nP����>���HZ�zG�"��;�^��5e�'5�QJ�ʪA�(�������r�[�����k�Q �ƍ�`��>�Q��M��\��5��-[~j������b�Z;��1Sd�F@f*܀���M��c�r��ì����jr\�����3�Pl��XTP�ru��?���C�,�s���-��xǬ0�/O���c�?
O���SV�A���T��M���{ �0��O:"u��MJկ ��S�/J���'�n����9W�N��F@<z9<}�����tY����A�A�5��є:���}�` &�C(���/�=��Xt�Зj��fj_��zs>RQsʷ��'�-'�R��c���
�� /��H�O�kmp=�6�e 	��A�.	�a]��-ziS�+]�Π�l}Xx�P�V`h�TXfEj����v��A�5Xf!������e]r̘I(�o��;��,�w|/#�Y�X�O&l�3���jk��Ql��S�P>��w�V�R>���E���턝�"h�)ݐt��g�D뵿�V�L����`���Ȟ�4d���WB�1�#�	zrA�z�R�tI��e!�)a���`�fűL�� 6�L'�]��<6��?,o��;K�j�7?����O#��V��Lc(0=�����3��,����S~hP�C���@�|���|�e��z�u�Y�G���'��h�E�������[�����v��xI$`�qF��Ȩf�,����a��eĞ]O�ն ,w�EK��m�5'��,0�{� �g�%b��bz=��/���b��K�`�^2�nE��N�m�J~�Q�E���(6�����,��"�D�ܓ���06���o���O:�k��4ʷxO�#?��-�jc
y.x�B���4Y@Ot痠�i���hƩsj�/�
b��]�i�F)�v�����b�Q5�����_��:��6�sKrl�JgO��,�G+�N��
�Vd�I�D {�]̑����K��e,�eX�J��f���	���U�y'�Q��ߠ�&�3�ܹ��'_0h�p¿Ι�|��[���$��7#Hq��6N�.ckտPA�XH24M=���8�?\�Y���b�3m����{T�qS�a����+�HѠ�&�M��߉���� �/� ��X�.2c�%A��h�k_�ገ��-��^�7��R��/Hߥ���>�_pQ��5��.�����%�l	���H�*��;j��'��PD�"Xa2c�{Rsڻ툊ĩ��4�,���p�#�k�����,D���&x�9~���뒯>*`, �ZYTFƨ/���M��AZ�MD���9ٍ�X'P.S �?��Շ�oSfNe��4E�y[��@܅�Le�	�[5~]E�hw`�x�g�~���7���jSFԢ�K�A�$ν��9mXA���܋y�3�]��7?����5q�Oȼ�7� 3`�Հ�N��M���Լ*�P�-S����u�r���W�v-:ӷ��dq׃�A2��p\��6
�q#��׏�=�z��#�%���g״���*	v�j�8�(:l��_�7�<m5'�˸�$�N�ŗ4��i���T���b���G���/K@���nR��#�6�������z�wos���VXꏿ4����0L�[a���?�J��8HL�	u���qBƵy�����u�\u����
�q�ُ���dW�a��:��aki�"�5$��!�E(��gB�Y��*of�O\��^�4��E���BP�6����(���}�pT�=XQP�U:ص[ ��j�-��k�l�ɼ0��H$p!���v�:�`e������@q��P;��`Fy�O_6w��l����+�I�Z���YĘ����,	���u�il(R���<ѱh<�᧡Q�^I�w0��vu;���R���3���7حl,����O2�ɻ�1+�μ��n�`\ˋ��o��1(�P��:C�R�-B�;��K:��|;��]1oq�\V���V߁)�\�Y���(��V���5c=�R�h@�&�M9DA#����t)����I���@k�̓gfj�+t���\���އ�;(]?��F����D�1�U�X���U
g,��Xo��c�����XR���g�-���ѝ��2n��l�MԼ�+7��&����Tf�e̺�Q�e(��}���7��"�V�6�n�HŅ�p����YX6?$�K��3M����g��J@)�7��������cq�]�N�w]�r(�{�S����Z)B�����4J�f^4�Z�7W�J�]t�!բ^?W�N�S� o�C#!�59�q�H�g�L鷸�/|�������v'���M�>0� 
	ĵYrNh�}��+1�`���k�Ƃ������\5K�L�~�ˑѧ�{����Wӫ"��	�XE���,ob�vt�����#��u�D�V]�y�׽��vK z����D%kI��iJ����q�g�'�Z-��8�ݠ�7E��ŭ���<Hn-�$ׯ���1���5tp[����#�� 5zu/u������2��4v�������0�!�����o�|��}�v��w-^΁�$�+�ϹX�ZÂ�8�dC�|ߋ�?8�5	�^\JR�M^�LI��f����9D�n�k\V��o0��B�Rh�c6E�
w1��2�AL���%�M;�� *��N5�Y(��R����Eq��K9�^�Ƹg�����Č��I�w�4�M�dW�Jټ�L������?I$��Yr�r����grN��3� u���t�����ts4��p�J՝�b�7�z�"�`W�g8��X�k䮿��0#_l�-��vI���8l�� <�5�A�:�����(�ja����= /v9��ڽ��m9�XV�O~���>v�~�lF%��p����J��W�ؖՓÒ���Z�Z��>��(K 	�$ie�C��:k7�d��ߍU�^^�u�/��ɧl-�A�]6|�-�H�a�iY�ַ��&t�E��{'CV3-�	W1d���\�!�.xXqw�X���b�pe��=�n$� ��҅ և*��iCJ_�[��ǧ�[\N����W��� �f��v?$��٩�[�e�N�G��D�"��1;Wl���z�����,���1h�E�(��Ô��� Dca�O�<�yd�(M��|wۤ�; gl�T���*�6��<��DP��D�_�0p� Ȼ���{
Z�u�M��֑�[G^TA���H��D!8��9��/�9��6��Y��>��V�����>��&�qǦ�<uQ�Щm��4����Hm_)�\!�4�a��*�^��g�=x��<�����M՞�=\5�Յ�Z�0Y�_���G Цv糞��C@��d�s`&c�ib'�h�Ro�^6��L��H]�?�gtܯ956��'�����������۬����%��,�h ��sGm�0�A�a]')�#V#j�{c����%�t]>��+�B�g:��[��9�h5�표;��9u��	ֿ7�m����N1�H�%�q��?�2vgNP�+=����Q�
��;g�����C�ܒ�+<�q�H�=@h���E�~�=pk���C�ݾ�E����QŁ}ת^�!��T�-�G����{0/>0�RAS�˩� ��Nz]f-uq����*ϒz��x@c�UD�MZ��O��j���`.b��^	��.�����m8���n�'aVҋ���a��ҋ����[����#t �'�,�~h��s#+us��O�4~`��.6o��NO�րpb��}M�U#j��-�ݸ����Z�t�-p�����\H��]{Kd�x�K~��7gMn	�7Ș�B�75�H���R'"��������ġ�t�-�N�B�1ڸ_s��9����ط��0Q|j�pۜ�%Z���;�ad]p��c?�⤵p �G̑MDӒZoiWx�J�'\kd���$3��*o�ԇJ�I���CG�57���a�f��{����[�YyZ�h��+�+.�u.�G��<��l7G ռ�������ɀ|+�<��f�5���>i\,9-�E��cF?��yVI����V�l�� ,�GX���\9�\���s�1�;sۅ��?a�1�ү)m�\�i|q;@�����0�;d��<���%E-������z�rJ*]��	����q�K;�˷e]�/�+/:�)v��وC9�ņD�:�#~��_��bEI���PAʓ�����T߽����E��:�8$5J��l��_EXCpf�
V��_�In�ß�_��m��oLi���!�*M�.�?����ԅ�K;��b�o����e���1�ɤ�U��fI�̝"z�Yfc)|��U����E��Q�u4j���S\I��y���ė�֧P�#1�A�>�ɦF��-�7&u�?P�$���:6�壒���b��J {g��ocmv͛��u]�����/Z������K�A[�}���NR�{%�?"0^�D�N�7B�����*��@�F�ª݉աB�kd?S��y���N*|nC���j*�U�*���a2x �2�0��|�&���T�Ah��w�����	1�w	���[�<#�^P��Z���z�6W��d�E�i�71��9T��<!��a�Ne�����>*�Q؀�#)�T��kPKDm��,m���L�v(E�=�_�9���{F��I�#�1�y�� �3~?U�	�ݔ�����^۷Զ�5�SE���@Yn���W�t���!�H4ð�%�&r�~v�(�<�]�ͱ�6��r�ꬲ�F���/K~�g,���P�~����d��x�t&���)�Uy�[SpLq3�A�Z�R�/��0�o0�/�t�Y���g����l�r��s�;�8������M�*�[\����;�Tz�j7��&ݳ��9XwU�+�h#j�Q���+��e	�p�$M�p��x�J<(t�g�K.۫l���g�6��̼e�;,eZ�z��j�cxq�t��⛜�X �H������$X����^ ���˚��o0!�K�Z����F{HeEnF�j5��D�4��?�Q���U)ؽ'F�`�r3��=R�kd�i����H�G&����u"��_��L숏���>��ټ�r��#2�R|C��ou�7UI�̵�=W��*"�փx�5{�r�kХ���[�;?޼>@�O6��I� K�0ӂ���fd4���Ǯ,��L��,�1ݤ/u�%^�v˂%yT�dv��)��A�q�t��I������C�nA�e�g���B#�z���[��D/�.E^wѺв"�I�	�%
�*-h���yZ�Ƴra���2���y3����]�s��;�Yl�����dm5�h�-�+��O�~�ܦ�"!a�Y����h�?�q\f���:(2>��B���6	���خe�[_��,����*��3��M�(�����U��Y�K����4Y�VA�_���������xn�Sf�R���%�d�jj��n��6'��u\ZQp���j�C}�/Ma.��-j�<?�oem��S�o��ݰ샣�ĭ�%�H2��H�m����_m��!�>0V���v��PT@��
0�=��V-���cp y]'���Z��6/ Q�B8�>1 �� ������J�q����C�c�b���Ӧ8���Gi�\�N��5w�=��q5k+Ω||�=�`��3�zg-Mqv4��ʝ��c//�[w�@�L�2��1�Ј
ǒ4�=�$̲�[��.�iZ+�Eo>l���FE�����= �8r����U�_X���?`Eh�:GK$�Ń�u���#z�Ju��͜��bt�!�O��TӜN���w�F��[�#Y<���#�/;:"3���D�����A��|A%_�AN"}I_C�\gz5��򭜃M]���0�l��������$5\�a=A��R���h���5�Q'�'x+�%�ɵ&���l�v��!��8O$�&����	y���.��r�3Un����21l67��6�,�v ��-H1Kr}�5\��c��t����e��X��r��г�K�R������������-A�N
�a�z��
�r�2%3�BS*���_f(E�'{&dn@�?#���:#!��IM�R���u8�7�S���
_� �5��<u�H�f�t�H�;��}
��֗ȝ�)s\�� ��L`V�ؽ�n���S�U|WNQý*�dwD(���ʤ*1����.�"TO���qg���J�����_Nt"2�u��e��c�WQ0��.hW�n�e��'y1	�-L���h��P>H�xd[o���93�\��
l�3 dG9�Ԟ�+����o:Ud�O);��T�N�1ʡ\B߂G����4Q3$�rC�=9�����Box���R���-�sn1R���<a2AL�L���j��c�Ʈ�d�O+㎟^~l�T��p(]A��1 �>f�U `nگｇ�j�D�e3�٧�A�3տ]%��e�X+\[S.��Q���H;�۴�? ��C�e��x ���3[?8�����p�6��b@�(g�N��j?��|��m_+#G.��;.m��z���e��X`I��4l��n��ňړ1FzOa��M�ǯ{�+ܸs���,�4˺!9�7m�6B�����V˅ߘL㇬w���$�!N��jn�'�\�\w�@��h�h^ɥ����.B��1E������Z#�hp��k�ŉ���(�/v҃�:�X�ł�:a��o�ö� �5�7��E�{�WR��0��aA������ֽ���r��NY��������r�5�~'t��Z3�I��U����Sih��!�q]+|��<���Jd�h+���k��}�Tc�3�2X�4Mb{E�-���r�a�;;m���5�2�v�?]�,�<�Y��J\���"��ߊ�ٻ�A�E����o�77�6���e��n�e�*���v[��Nr�H�^����M�(��q�:�W��S�8����TU����7�f3b�u�d�X�s]K�&a������'Օ��V�a ����uK�@\�NG]e}��*O<g�~�咴��X��0f��<���w�D���#C��Km���N52���"1L���Zc�ɿq�����(Dޮ��5/H( _� �����5SLUyM�K���E�3�V�r�$�*�'�OP�;�I�jP���oE��F��
9��T%9�{�8-,L�I���]T��.	�Z#am��_I�m�o?d���XV�Z,β�&���UZ��u-`r���++���3�摻*_����7&�<����	e�.��M�a�nt�������Y�f��;�\^Kj� �Q��ǕL�|M]��^�<�D����*@Q�=����������<��9�t7�xh��!oҹ�,�@�����Y�iw_�K�z�J!�qL��SOPř��d{�*��r������g$:	%"P�}������4��8��F w�D^^O�� ����o���15>�ne�ԧ�$�`z�f�i�\�[���e���i=���r��}M����C��ڧe�[W͍ols��{:�N�`g�l�D�%�T�8� 	�j J�0My��s����U�
����Nu��N>��*2�'}����e�1�r�����G�����DFpb�{t������]
$����o���2a�ri�6�O�F�x3��IW "��n�!���^����nb�� e��G������Veu���'�wT"`�ۇ�&��cdt��a�OR��³���Z�N�Qb~.��Y#f�K��
*��(Vy�e3�&��E��8D�u���0p^`֡��WE����6>\ݤ� ����}�~�ͼ!p�cd���]t��L>7{�x��c�m3m����M
y������H.*�����>ч!�Yr����.�%WQ�Y�{�<�ƛDd�[�.oc�b݉{��9��_GX�jj�kJ�t��M��U9���ѐ?���[!�A��Zj�pj��X&Ũ;��x��L��G*��3��8�7�����D��"7VF6���:
Х����M��j�kw��>�!0�R.SQW��l���BY� ��щr�������Vl�/f�O��.)�	�Ng(7|T��q0z�/�o��s�U�/Q<5�8�ῆɕ!�_ ����3���Q�B�N�0��i�VB�*�]��C�([��u#<��'V&!��?�I�AJ Q�o�q8��9��eP�����V�����VV7)�����:�ӸaW�캞ώ���	�N��ed��Q:��zȯ�9�0��=?��>ɗ�kuw?�s�4�?'b���)��zdޏ^G\]#��6���ĺ�ˆ �^����]��:�L��g��L��H����_*gU0��kK��"6F%��V,�,�9�/L(/,#=�4����֎}x<07��p��B������������x��؃���{��a�y��O>½��Qb� i;���<a*ή�\���9{�A;���,���_k1��/Nh�ՊT�cOEB8�Ѕ��Ua[m�]T�P˙$�Y��Ƅ��^���o^E-��7-����:j�=�~����~o�1�]����/҉ZB���_Wp=�N�UQĸr?��!��.�v@�̪fc����1�(V�:L�rbZ��H�o?�@ D���R�:���<dJ�C�QAҹ���+���;�����3�H�_����<�;�څ��4����[5��:��r2?W$h����>�;�a�J�g�VB�� �_Jû͒"�S��mx�!�,r���8�;Pd�b�x��r�JV�ё�gO�ǧJ_u;γ� �M���EÖ9 x`N1C�rN��*�$��<c�������1�/ǜ�mɏ9.JL�`�ue3�N�h�hx��3����8~�)
�@Dnƻ p
#DV4�����n��tޣRr@����xN�@�2?<�Dd��cu�0N�Q�&ç�Q�0�͐N䤇j�8v��)�U�C1�>\�Xfu~�{���<A%��Y�x��	�3�՜׌����@������>.����
�m9~!�YJv�:-�uf�s~�� H�Ό��^k*�u|�s���p����<��M�5�Ҳ�N몘��T���@{���şt	�c:�kL�%�o��\P��+�8�DS9���
����E�[�U���o'1M�\	��f��GkG����T�WᱍD�i��4�o�&���ŝ-^,�9�!��N0������F,a�˭��?_���mm���['���v�͖A�-c���fr�7��~| ��ӏΙצ���.�i�Nb�r1���.~�u�ɵU���io�8���p����<C5����ApBi�!��*������;k<�9�OrD^�R��D��6��}Q�P�("(ԏ�O�Ċ�kfx���]��$��V�A=��<�}p�%�o�X oi���B�=5P���z!���1�{����cE4���U��!���ఇ��[�9�1��I�b[�;H''�N3fO�9�\�g��f]P��84:c54��g3��
Z9��D��,����kO?�]��TVaH� ��(b�� �ư�U�	n~�X�I5/-��Q+�I;��TE�e��o]X̏6TW'�w8x;b����W�9���߾Q�t�{,���kмC5�D1Y�L�D���J��J"]�N\�0ʙ�G7���I�y�PpE�pS����,H-�"�W�f/���ņ��<=�J��Yn�Q�,�WBf��8���E�_
�l��,��Q���3QKRw�c�(�tl-f�!�ؤ�]�U��ϔ1ՍA4��vޠ���������|��3������1>j��h.8;� )�J3�T�A���8W����{
�@ �%��
��%���Cڼ�`a��!��G or��ml}�y���H۫�mf�/i0M5~ O���$����"��a>��ʆT���.�Re���o&ć�`�+��;�keGf>i�7;�����x�Md�X�w�&P�e|�"H$�炠H{nƢ쫂/5�5�;>'��c�����8f�&�?���؃]v��z>�֏gF�h�u~������9�i�yT�]	�v1���3<W��F�p��?C+��u:��#�[g��~�M'�<\���Y��%�� r�����HW�,t6�F��xsh�&��U���nCl�]�������7��i�U�E��<b� ے@��q)����rK[wnC2�9v^�i�H��))%Q���2�H .�*!��<"�E)�J��n�.0���83-sb�W_�a�B����b��_>u������=ؚ�մ7�[�b<f ���8
ǡ8@��)ƻ��'�Σ��A[L�b �Qm�2 �!e����c_�"�a�i�,�$Tb�[��_V�kk
Iz�uB)�"S1H�}�^Y��?oF�����0��*��YO��x�\�d��%'˒�M�����(a��A�P��T�a�\��;MKǥ��y3kG��>�����ɪ��q?9�����B���$�b}�?E<齌2,�Q�<P��n]��0��HH_��Lk���m�f�>x����w=���?]�q��|�(r��,88V�u�O`Ǿ[�*��6A?�_��G}SQ
�J�@��#�=��y��dA@{ۋ��b����Ǵ2&���8c��f�1f��A6	?A���t�S���D���~�4�g��8&��X��:���x_��[މ�+�Dx)���\����l���	D�J441���D �&����&���|-��Ӯvwdۘ`'"��K�17G2b��g��
�MSIk�{��pIzh\K��W�����m�ěW�S)�EGM_�0��?9	�n�V�U��*��ȀF��u{P>/=���5="�����C*�/�m-!�:�f1�C��3f)J��y�JD��p.$���K��xΓ𼙳��v$�����l�.@=Yl�yF�s���bm�T�	�A%3ʉJ�n_�LzI�{��Fiht�$!��V.��+x�,(�s���=:��&'���(.��ā�Ό A�4{�h�����&�rNP�]j���M��^s^�`AV-V��]A�>h�	rR��.|֊@��g?� �+�&�orbG��+�i���iMAo9�i�j�z	���:��6±�|�Y*�o]��ʩpAcȪ��ag��J�xUA�E	M�{�3д��������K����݄�O����h��.$D�{��[�(�&TC�D�վ�>y9�4�7!��A9���Nq硔��rzיM�G��۲�g;�lB��z��mc��g���sm���t����={�ZI�T��C���LV���h[�1�E�כDϾ��g�h�+�ĕ8p�1�5��ݖ��0�l�d�2��>�x�sD ��������;�)�X���}�(�?c�3���mٺYk�3�M��VL�_��Q+)��~Z[�$h�+Li�ǙB�n��3���?��f�~JW�g$.Z��O��������/��@I\�t[t�6�->�sB�6dd%�,��4�TƳ.��L���.q��n�~��Z�����e���d�BHb��'p�[k4\��(\ܳk�A!QJ�Rj3�Cڔ���Z��Zb]
�.X9����O�9��3c���qJL|�hZE�u�捑pyb�}���y�!�I��0��1<�=�W�u<�P�5Ԍ�;�g�y�jT�@ܜ��僑��
�:��Ql)K-P���� |�H�H?��F�g��k����J�~��	~����;�vf������u�j�ߍ�UO���M�pQ �z�m�Y2��=w(E� $+UuU��C�茢q{�#	�Á�����z� ml��.��7܌��M�d�3F��-t;�$G6�pѓ!(���pwT�oO��r.��%�p/��/��J[�ţs�s���H�U�ޟ\� E��u�� �p6Z]
"Hk�#�;��T$#M�����`7 ���3}`#w?9��L����fhۼ����}�卉���]Ҏg�Y^�M��g����H���o$���5�!�����i����b��Z V��U�0�b�`� X�+ ��]���
�h7� �쟈�'QWL�q����mK�j=��򚙀���(Sl��w�\��׷�p?�E�2r��IV1W��w�|������hǡ��B�Gy{�������a=yx���XN��SM�����F��)��[�~J9b`nYE�1~����u��;�=_�A;���yw����җp�Zv������N���]�&��Upa�����#�g���8<*�u���z$.��3�9�͔�:�v'�����	�З@�����*�+Y�A�ֲ:á�Z�8��o+�mì����LbG�f	۬�U�JR�p�4;�D��-i�3��wn�L�9^�zT&��l�	�w���4&q����������NN/h/��ZY�g�,����za����iby�������P1��z� �ͱ�.��)6�+#�/�x0~��6rʊ"�,El�K��:ki7�T�+�l�.�҄̏I�	%��^����}���6şt���D�f��Y�L��5�EFpr��`˄��qH}.�ٷ/bٴl�Ln?4NH������ƅ&�\=F�A�����L�ur���y�]��*�@Ӂ\:2��F��v��y>�jf��MN��������]]�6+͐��'.���DE�Q���V�4:[�u��q-
��;��
����:|�"���;?7��<��]B�Rҕ��ZU�B�z:�������ݚȒ�м�����/	s��N���߽����*��E&���ؐ���%9�!
��VȮ�n���΁��r�Ak�1�����
�zqi� ��-�i�G�����O��9g�#c�9~_3��<�F�s3����h;)�R?��"cܴ>���%�`�>�	Ѕ.<�O$�w���i�>�Łf�fF�Ks��L87QK�Q2��}{�4lZꮎ���	?�g ���C	������\KO��$�
/4��< ����q�V�)bL����l\èpt�	�G��mn��L$ǰg����/�p(�/Vz�T������c	�O�K��ե'K�C����`~��y�w7Q#�#��x]��=~�
�3䣤�(Evv�����%�j.��C��{H4/<�����W�P��5W�9E5c�t�rX�`�T�̹��:U�UZ\�dPx~��m8���:���k,esP��b���d^v�[2�iZW H�`�шN[��M2��'-�W/�A8�qD/��׋Ѿ*q�k���O7|H8��2���SRT�0MFݥE'Yu�7ڬ�,�S��2��/M���8��+�^�o/����	�;�I}l%��g�h��m�e�g��ԕ���uX:/8o�b�Ig�^J�W�aG��V�QMqO!*(4T��g�=�Ɋ����Q�ƞ.������$ϛ�6�C����c�x�A*z�]����X��{��;+�6V�P	l�;Y�//�U�{!i�톝P�H�δ\T�`�aߒ�،������t�]��1c������V��/��DL���^�	@�=IH�E�����9*���0';�]�<(�0��E�j8�PB,�֐q�`�h�0F*��؊�.��A˰!��s"�2�r�jW6���G�xD����_�.��$"Rr
��خh�������}�:�p6�����c�S�s֌�~�m#�<�l#q�"�-ٕ��8Zy���y�j�5*�B��,��(�Mq���ppt���|t�\6*�7�P��Vzr�Ŀ�!�%��~�Ias��6�=KdP��Q��Q~`w\[+Q ����%��I���H�������\�	A�g����pZR�	�x�}�|����"�}m"����A�-��(�(U*���I�oI���؎�8-�i�(`��	�;V�d5�*���� ���	��k¼lօY�eK̡�Ey�y����\h7�c��W�Zːޛ�F|�L���~�_&pQ`�����8�K�%{���kFn>�H3ǭ�f����5�/�(:�"#�����j�\ғ��%��!���m�r���"<|f�=�ܝ�u�@kBB6Ss�-T�XB0�w���;DO�dc�bV�QV�
�י�'-�9���w�҅��X10[��  ^Vb���0ն(�S����~�T:9����w/]5ګyd5�۹T*��ٔ��R����H~E[n~��\���sg���p��+�)�=��L� �q"��M?��\�6,7��y���;�/X��Xm��J�:2���i�  ��tC�3�'=��V|�#i4�/�#wJ�mS����籩(��cK�o.�D��u+�`?� **/l9��Z|`p�6�����*[nȹ�|9p��Z�u���a��^��nw���߯�O`$Ѭ��[5��3�U��B��k2���A����`�i�(�$|XÄ�3��Yw�
���mvg�x}�/�1�m���
2m ��ڶF�����x�Z���1�avӖ<���XY���|.vid|�O� �m�0�e�{_mp�s�@gc'3��{2����j��#1�s�x���-Y�$�FS��Je�۴�"���*@�y���8P���Fg��}�F?��V�h�Ke��4'��r���� ��z�8���-�!��6C�s��%��z��'e6d��g��s��%^�G��V�Ë2�T��d�<z��<�䡮�J�pz��	P��z�
�z��R���`Ϻ�o��Q�vXP�am� 'ľ{����/)ԛA �tn�3Ώ�U��8��l�O)�-F�<l:�ۮ-;5 �ю�,{~���)�*n�`[����W<�_|���:��g1eCE/��Y�=s��Y$��yd�=��v/ܴr��ju���Hi�֏�W���n~�����1aI�����$s�M�`��R_x��2ˣ�O������{~1�ީH~�;�Z^�t3s��Ȳ��43�e���@d���� �J�l�X��݋z5�G�W0�PjU��y��U&�� �s��2���6�yB�G���ކ`E�4Ӹ+����w�ZQ���$������E��_Y�3-u�@b6�O��t���s����y<��ʫb��ujx;�t;��r�kHL͔/R����~(�xt]��f"�U���ZNF�Ą� ���V�3�6=$}����H�,e��W�"�X��T]���,��m{�a�B����hȓ6zI�rP�da��z����Ql#a�EX�=���[��iىH����1s�Y�ŋ4@`0q�<��&�d�<���~+!ғb4�B��	��Œ�ej�Ĥ}���'�Qt��jz���g )�%�S���4��v���w�y7.ҿB+�Y��d����h�d �� Z�L��"b��N��c7����ո\�<Ӹ٣21P�,����e���*3o�i��-B�?�*�Uf���mzmq/��},=i�����5lw��ǅ_��rHfM�,�?LWW)^v���b�i�ڧ���P�41�� S��uq|Q�},@�;������g�P2ę��B��n����Uύ��I�f��2i���3������82��R\y���ϕ�K���\o��9]Zg��� ��GUX�ȇ�t_*@�3�mA]�{���;x
��PQ���F��uwTv�\�u�.2l@c�1!bO�z�������2��:J����4�r�(�����K�H��[��7o# �j�.Ԇ�Ի͌��{Ċ5I�l��^�B{Gw�G �Fo�`���=`���ɘqv�i��K���_�8%@���SM(�p*,�<���0ڀLl|2gt�$ߘ/Mٽ�csn���ǑqM��1>�8��w�S�r9E��#}U�h�����_��Z�9>�tA��`���U��&L�8����r�C��Ts���Oi��Z+� ����&���G��N�<�omfh�:�X�0�x,.��ޘ�F�Zc� 嫭v�G4��.��U�v��>~�(`�y�y]�?�~�=��l+�NFB��QZ�#�q��Oz��.D��Okw��Z�7q�q��!��הPZ�	κy!�<z�����:��7��Z��Yn���/��A䜤`"WH�'�����Z��հ���%�t�- �$����l/���;:M�Q�r���ܜ�k?)����,II2g3��I��l�a׬���'k̯����	�2JCZ�(Jz����9�b~�fc��= o�`a�� ���UZdT�h5��� ��[�R~ΟW:��u�x��>&�7��>��v�M/�6���xPA�Sc]��G(���1v?�#Lvf���-��Ǒ���)d!�kHO1��vL�!_�<�u厝�۴���Y`���i�6�߀����+�Q�z>��O��ᢸ@
��(��X�a�Lvt-�`��������4U�Ȑ~+V����]��>�����1.O~-��a1���r����eZDp%7�b��||��s�OoF�`��0%�e$B���4���[�m.<���iθ�H#��K�̧C��2f�D���(�U�����G��v7�P<���iT�� _����&�d��_����%��ߵϔ�*O��H�8�ݢ�V�SL��x&���)-R�<�5D�X�9�y���Eá�
�H[�Ɨ��y��ɖ������4�	y��;�ե�Ē{;Ҁ�#�D�����VV��8�B�����Reó�t1�.��aQt�&��@��c�6T��q����������N�E�;Nx�K���(P�E�q(�j��g���|��i���qڔPxD,j>-�auB�����gP�����\�c�f��AT�������vj��)W�o^+�%��7�{-~"���P�/�2,�9�-�fy�*}.#�KL�A%�X���=�Z0�%A��(�t��=��n��h�6������8�mS-��a(�k����Z��>A�x�6�����+��#;tָ _����#E��c�uqcF[�ms?|];LA�}��8�sG��K�������������D�H�07d�;��cS��~O<_
�a�i�n�QV�0�]#�
��4^��Vvok""�gB[*�o�Z$�8�+��%D؟ȳ�5��nt�F�%��� ʋ��ޕ/k~?�뭓]y̶�|�ųL�B����C�9��6�����u�T|O��J����ԑ9o*��~�j�Mr�m
>}���)�c�YȀ�m�L�Q�F3̤�2����͡?@��MNA�R
(��j|����DB� �r/�V������b��o�z�������";�%\?5T�����ء�4�2���oC������kjʕ��~��0���n�mҖ��~x�{�}㢤=X�x9A�����Q��w�$Yw�Ոo�Kk��	����w�A��6�7f�w�G��7�/KQ�o�I��Ҹ��J��t�1���m����I�WmV�Y��fk_{z�r;{���Η焟��w9	DM:V ����㵘�ˤ_O�7q��̊�w�n�{A������i8������
�q��y�#��"\r2�����\�vɛ�$��2�G�%�����P����HPM��d���{�e)O��\w��^S[��3�����#�Q{�rM�-V�Q�b�van�=�°�Q,����t��Q�&�� �Y�i�����$�GïZ������L`y�I{E���tם@�.�V0J���᫩;^;�Y�š'�O�Ay
[e��/Je��of�r�"ѧ����0�+�#�\Py����I�a��{#qp��r�qvE�ysN��s�Uu�byYv.�D��!�R쿎�� �Xb��^���[�v8�(g�5�D���3-�-��kf_���|��h卖δL�|,���pݧ�O��"��q`��Zg8|f'id�~�;r�v�c�M��/*����bw:�נ��uW�I�"SwL�� ���gE>��7o>���E��9����ɛǶ�-tKD�N>����i��~�d��y#M���Ll�J�M��� ��c	c�4�u���=5!�gG]��KG���]|f�]�.��DĘ}����-�E_�����P�"l���p�p���-�_��g/d=+y��D䷢�̪��jؤWEBVw�Yα��)_���ImFz�~<��� �����e�J2s�{j��gI�p8�ٻw���L5c�{|�nF'�q������ﳛ��kN���B��e��]c1��"]f ���%��G��>*���F�M|��C)[�=a� `�����S�?$fj�dص}�|ls݁#�F��� l9�xL�!������*t�R�77�~h:�&Ar3���=j��G$�@�Ó.�[jM7g2	`"0����dxZ������̵gOD��3~��o��k1�QJ�����}V�1��ۗ��^�:"�'��ō�y���i �B�ǿTș⭰'���$������n4 ���F�������n���_�9����-U�jb��c�<�7Q�6� ybV��q�3���ʸ�I�,?�ѹ
ڣ�+�:��TZE@K�o���~�-�v���l�s?GV/�9�_0��@�+��b���Z��W��2�'��n�P
F�ʔ��O�֧��#9�U�܇��(���^ /�{v1�w���Q �$��4��:�1�Dz��=�^��f@�e�"�T�TQ�d�PC&C�~_r���ͩ�E�)�6ڋi�qXF��G�xI,�6m�� ��a��<�����4}�	���hS���b4����;�;�H�:�[���&�+�!�f揓q��e9F��,K�tk�T�M��8)���h:�\�ל�UӜ��9�U���T-��a��Q������=.�n2Sg����\�u!V^X�g�p��j��i"�cF�q������\���Ӝ���	��'^�oW&�4>�tW9!?��%�b�>�9�L|�3��b�h}_� �����,�
�j
E�Ö��6����=���H�tj_�k���S�>���#���*6���3�����"�s�G����r>�?<{.���v=5��g���ȭ����)L m>Z����Fa�Ƕc�C�^p�?�F�(.�zi��Å��`��b�\�4�QX���vt�>q��z!u]Hb8�v�F#3�h�t~���+8P��mg]W$Td���C��Q�� ���)���+	0Ќ��~��U�'FkZء�����[gB^j���������,ؑH�2���no�����f��׏��E-�Y�`��I&��O������\^�AT��J&��L�d�	�ڬy68௕w��г����'��#4��d}��ҫ��.�����ǥU�T�t�x������(��y��w�&,aO&�3�E�f�Oy��S��+�[OB�Փ��nw��cܕL���y?�1�%�q�9�x׸��T���볛nլ���q����O�k oSB������2f�yH��������|**6��\�`-{�`�wvu��~�ef�b��z^h�����	6h2K}%���+�r�� )jIF�b�	BӰ ;�{n��̷eZ�<[p�`;����5���ijh�YRf��Z���<�uC�������lL�A/Z�,�)o@�<���i�d��`J���&m>���P�+U�.��:>S�L (�-��ۿ���*�n-�V��n���jΊ��v�=�/2����h�xbX�á{\�z�:gUf�
u�V�y_�v/�M������Gns0��+��)]׏�)fm�-�a����v�XG�?�Qy rC5`Ř֡��������Z�/�6�����LH�1�/t|���.�i��]D����]����P{�<�p�5�D��
T��$1ku��).����3fT��8&ʨW�`���(B��Z��b!Ȟ��X�߾�L+8��{
>e�!�[��E�N�S��I`e��z��tW��a��X���Ջ�l���_��e����$"��>��3-5f�Ě����%'������I
���࿚!�c���/Q��q[��6�e 3��C3X��:��9ۈ�������mM�A�<�Z/�H&�`�xH*�=�����7��Z�-{��(�,+ؗ��l�6���D�BaLr�દ]�s�B���P.����8���N��`�C@����EbuI�z'YdΓ��Q�^h�w��,�O
L#p_*K�c����G��(�*7������s���޴�������X�:�^�����Q�2�]�/|��� ���v��E�nX�-���%	�:'�#�FN9<-� �']�F��k�CpQ���U|tUX-
��,Z��7Z�&Y�j�T���]hñ����c��`X���tk��=1����Ee�C@��?ۘ��ݞ���
������k��ZD�w���P�8
Ͻ�^&�rL)� @1٨�2ٵ�ױ$R� �e0�K�S��&�>�=_K�W���b�d�ء󭰱T�?	6�F�4�^���!C�ɕ~�z�k_-2�K��Z�K�+1���
��}X3� ֡��^�v<�q6�5<K>�7٫�}*";���~,�#�묽EF�]KtrU��(� 4��ʂ��`jF'L��@�ɬ�^2���݀�����<�k�Jξ��V<}Y�k�>�:�T��G��������G=4�bL��M$ʹ�l�N�߻��l�J{:t�s��E���p9�R�#9�u�������юRԤa���&��V8����|ow6z��˕�`�& K��rތb�Z���	i�ϫ<r{�,�Y5Ӭ�9�yBS�k�qW��S�ЫWӉ(E��|yN���V5f�*�o&��Z�09.d)�_
xGb�>ob`�]��]N��j�-{�W3��4���#�{�j�V��0M�'#�1t��NE��@l���{��Z��MNI�ܻ��DϾ��n��ɸp�"1��:�#�|����
�:{W0qw�p � �^p��w�-w����{�}2��0��+��x2��C�lpv�A]wF%�S�	YֹV¤I�I3���P���������*)N�{�Hkx�8�l��=�e%#�Z�IK�<j�v�=�q��:Hl�����r�Ҭ)C����+_���ϔ�m���&����%nv�C5E��^q�ݲ��}��&f�T#�~�L�6��/�l1Bj%���D������/���D�Ν��_�N	��=�5M0�@r�R@I���Ú���bϼ{�.�|W�W��C��r��Џ��D"%Ǜg]v@��{��*�`C����b���0�7���������:�*��&�X��}Un�L\��0��4&V��#Hݰ����sh��e��&^�_�x["�Ih��3s��-ͦe=�г�gw������������Y�����*.=�6]d�=��x��-7��,ۊ�����Џ�ae�L�T�:	��AfCx��F	�k��UB�����v��E@�.��g�t�2q�sP��8;F&��}d���k��	��	�%��W�����:?"�,�g9�xGfNZ�
���t{F��@p�)h�EO�~p�䌵a����H˽�6��2�Q�;�b;B�0= %5ƌ��-��^�!�3>�aH�w�F��K$�^����/�(�����d���-�|��C��qg�ύ�,�C��fP��[	z�ٳII����i��ޚ��D|��u��e�e��z�ȧ����w�\��l)�{�B5q+��p�����:����D��U�i�:6:G�^��s���BR�������wN���).�1�g-r��I�ܘ_���ު���gu�'Փ���֨�V���X{(��`�TZ�Po�7Q�k	��_a��}��۲�0�)�ugzM5'q����Ŭ{�n�`�ʽ,
��/�v�`;��]��KXB&-�Ձ����<1�+U"cxК1�4�G�`�o������W����Zp跟k��w��6&7.��<�jd��tš�努`��&Q��U�"<��v�N�Y8M ��Y�����^��܉Jn]l�C7D�!�Zp)�ZA\�ۇ���q8�8C���6*�����%./*LɴX'4���"�y$W�S��w���՝�h�6�����c�&�m.Ni�ԯwLԷ�P*<�V��D3L�c{���v��q�̼�S�����칍�����ʓ�oW��J��(px��V��q�Ӡ�o����m�{�{�xQ��ᮢP��}��/�jʥK]}(L�yG<��o+��^7�id��8��h== S='� r�b��d�� Y�,e��V���,n�@���af(��������������L����q>�T�Y�ٛZ�S(��wI�9���d�JP6m"sC��"��^$�-8~�_f�ˊ���B�U�WO\l�|�x�qXi��eԔ��k!�R�ӉM��h����ٽ��ʂld�ԫ�eC�v M��`r�UL�M��.1=]��LHAdg&��D���oly�1��Z�<��D�
s?�lq�_�䩷�'>��V㮉Ycby�����zh�4�O
Yv��b��}W������e��C��5�n�?�)E	J+�f"��3�ɟ�ADß�6�Q�K���?�E��+;�f|�ŉ�v�j-N{���G{������ϵ���s|dV�	)���y#���:�P��Ս9�y�F��▹Zp6��� x�I��������Fh%�s#2_"�w�dP�(k�n
E��Ȝտ@���C�7�������`:Jo�E?^����]Cu'�|T��+��8?zx���H���v������A��UM���Z�&����2���gk��^���Lh�tjDA7F����A�PJo�_�cXj^��e%��U���/u�w���
� ��8C��niB!���2ۊ�@�?���L\IIT2t!��TYTq/�tK+���7M9���A�f�S���Ē.q�3�ـC2�^�mj�I>W:��
e��gc�������F��Y�W��G�g�t6g���fId@��P�6��(�Ck�<�;?�
��؎�,4���ͿC�d.o�N@�M6Ҋ�7��$d��Ztؿ�j	�K���g~�Z_і���Xի$�A�]�� ��YB[���FR|��F�:� C{�z�<8�um��k�Qv]�*����A���`2��~�W+��2�d;�ƍ$�s�!:�ד���C"�)�&8�� �w�,�`S{ ����N"���\�&B�.��@����MS2�U| �CVW��f�Q?F"�saY4�Qӣ$t�@,"1(�3�c���f�s�.6�D��B��y@DI���fR�Yӽ��Jqp0A��?�b��d\_�S^� '������R�5�<M�à"�bTJ.�<�E9v��w�1ƈ�Ef��W&!j����Px��=2����3�<(�H��z��x6�}��A�*�g60�*�����8a�J斒�dT�_]�'��}0�3�	�����&`�KYn��`�;��F��v8)[9j�����ԧv2� Bs��Nv~�\~�:-a)mH����f�H��[b�ry��Z�ح��H��]踗��)A�TI+�	��ɩ�n)��T  M�V�!Ԑ�KN����PǛ��²PG���E����jDj�$���,�\���íJ��u�p����7h�1�w��6w�!����=�6
�;t�{z\�d.WZ�?!<����U�߇�Cx�-��pm6!Z���J���.�,؍�~����(�dڽ[�C�Z�2�!�ŨPk�`D]��GIo1�(P�[2��vӊer��W��8\�
�龜�/4<��B�p���Pլ�}��]�RZ���{�#�������ݸ������r;�dL�W��A��h�N1�4��.R�r�:��m�+y���m/���
�4dӓn>��a�A�1�	K6�M2a$W^��ق;�j��4<{{�����]H@K5K��ٷ�1����כ�{?"ɮ�"� ��|8p58�D��B���&�'c��7�1
�]���h-��8�{/�ha�q�b�=���>�痗�(c-y;�]W)��	���2��M��H�ĂQ��"�9m���M��h�9	�ۃ0�v 4�@�-���8�p2� ��������z�:Q~����)��k߉�U�\w�}ŧi`I�cw�n=�>n�m�;z�Ww�>_s+�9�n��>�N����ἅ(��`Q�[C������Fl��v.��HI����ǜ���P>�[cd��C5g�&$��Ҕ�R:�@��z�1�ح�vع�������5���洖�:G!��Gs*3�7�`dQfe�'�̲C(5�����}�Z���1��,+Z����e'�?�nPs�e��b�?����M �PN�i�l���G��	u�̼��.��;�p��&J��D��41e�@��ճ%_�2~�*�3̃6��K����D^\�N+��� ��m�//\YRڝs�I�����4�����t����������K�l��D�V�
_�Y�� H;��!vGr~�Ƥ�ы&O�jBG��O�ϛ�&�Wp7zO1Dl�T��ȶ��V\�>�&4�%PO�
K��'�A`�Y��Zi�4b��RR�(#8��ұ�W!:'k��2�J���#
�㍽��#�W.C���NPx�@z�U�H�ٸ$�ƿtzF�X�`
]��K��Ggz��'�mZNn�sZL�9+��%j���w"y��\?� B�s	��ST]6*��^��H�U�Q�����Ά��l�qUؗӈx��F��������4��h��n�F�{p�l:�Ɉ�}:"�z�Ɨ�B늧�X�|P�j����s@X�'����M�O�&��j-yLؓ��0.��������B�S|x0��%g��阶�)g�kR����!N|wT(�3�:��76���˪@r�2"����yN����n����%����.LP�~(h"��֨��H�5c[K�fT�F������[�|v�XKU����ݕ��.OwY9lP��Ꙛ��ho��g�):p?��`�L���DvV"yB^P� 2Yq/Gs|aM2�,�*�Z����:po)�\B���t��pf�����f= u9Z�;Fz񴋤�
V�4���1�o���|)h��'�`<�9Z�zW��Yj@&&t�*��kf�X�x��w2ԗ)��n��2Z�0ջΎ����kɯ}�� íP�V"�?o��nv�~;1��ȱ�3��z�sЪ�RsU�Ĳ������oV�e�ئ*vU��?l�et�Z\4����_{515��压W�Mf�Š�bKE��)4����R�e���]=HPn}� �Z�aO^ �u_^`��s�M�)���<	P������6�+�� /q��Hf�ϋ��=X�O�����,�!�z��u�|�ډ���x�jf-Z�-~+E!y�q`%2�	�smR��H�]�ǂ�|��u�E�P?F�# �`��S���c�&�8)��ĄC��I�c���}�ԃ���%�7};8xW(NY��-Ż��e�����S���[�+����U6o�m�?����Kn��!�բ����ov�����9"v,��5��ߪ]H��/��c��1�=։�xU
e5+jh��9�%:�q7�m̛�}��s�z9T&�D>�$�#���*���3n�5Y7GxD���{z(�-�[{QU'B��a�aT��c�Ki>��4�QI�I5�Yk�F����T�9�s%��5�Q*z,�-<&|\	V{񡓝��)�S�7�h��WR��C;�+A���oO�f �g��U��OS������5�7v�2�.0�e�6t����/��;b�d�CC
��GyK��M�H4�]����t��$r�@���PaWr�ʄ �n
�ϳ�%o����~��^�j����dpL8n�&z�t�e�<�|��N�Lf�ӯ�������R�3,M�]u[W6x�L����q�"H4�`�ȩ�~��R��*��4�H>)���'�r1�/��{�!:�l�u�R�� z4Y�I'�����I�?!�Ļ���^���ӎG��I����r�������Xݞ��xg7��DK,��X`����r�r�aV}����b��T��@�˞<��R�8{.ػ�`��e(�6��.�<�Dg�ѳ�����'~նc������Dk��i���k( bT�1<4X��N�κrFm�tk��md/)������^��め��
��[(�Z�f��s"ѧ
^H-'c3�o����h'����^w/�߱����� g݉�.*?ժ�6:�y�w�fލH!�/fC_��fMuX��|ԻGF�[]�_��B[�|�,'�9Uh8� e�����Oϡ$� �P&D�w�`����w��&�ns��uLS�)�%I7����iط{�%oܵ͞?�O�����eW� -,�W	�:�fp���g������>I���B�8�SF�P{`;a�;n��b�������P��d$vO�Rm[ʠ\3�Ἅ��x|�ʹq��~wFO����7���;�$�� ��=`���``a
�B��nL�`
f��ߥ3��y\�5���5��.8��U�s�g��ʬq�������j�����C��_��B�3����9����ю^���4E�g��:���%��b&Á}F_��D,�q�#���i�7���x"��c�����/kߗWK��d���Z.9���'��44�$�'�ſ��b�	oQ$�X5j��P�ϩҼ��(p���m�a�#��f4��^���K���!��
S�s@aL|���}��sOTe\e�ـ��u��Km�og�H�������S�S��]��z_�g�1�yԆV��DKO2Hy�lq�\%�����H�pg"r��=�&�#�DEY��o���Z�FY��U�@�D��9�"$ ^�V��[�R�G�BnYoQ)1� �-,*�4!�9��:6��F0���9Fg��T+wV;=�9�������Z��߬4�!�vҾm�3���"��{����t��]�8L�ZaE�q��}�L��:)<�O�yGzW�a+�`�d	U�$~��rD�P@�"�K�+�A�ݹ��~�Y�Sr�If?�B��D�e���ol�%�G���70 ��o�]���}��8�G.�װ��_Ǧ[�h�+��U>����;��,C8��FQ��iD�dI �)1*�;K����Kw���_uŵ|����H��̻�"��~bx����<n$P��K���]�e�s�H}ڨ��ٴ��� ���a-�f"ʋ%���V�c.��8J(�P.�<��� ?ۓ$���2^���.�v�wt�M��O殖�Ϊ���F��τ�;#wSP��>�ْ����c;G�) �k3=3�:�)���C�Ja'wB��+n�h��o�r'눺�����z�m�����/�`����7�[,̦J#���}
jy�D���R�ϩ&[�`�/�C�0��?ʣŨН �穜�LC#a͇�h�H��z�S�X¥�o�$�>�$,��#�|i*7\ɛ�K�')�rf1����E	pon�^��K
�f�n��Rd~[�^��L5dwmz ��v�\�(����Q(50̺��o�y�z��G���z�a��-�r�;�\|�Ļh�]v�淿�P7�c�R�!)B�{�E)Є"��E܂���۫�y���_\�v�Fs��ܛ�E'(���K��dµ�lM�|E��v��b��r��
5��ݧ�A)�p|q�7��<��qxF;x�X��.�<�1��i��I�_)g�vEaB ��v���Ҿ�%�q���-I3����b�:�wZvx���X�G輏RY����gt�� �� �S[Ꞧ�����i�N9�$�ZR�-�����b*$!�,��*Ѳ��yqiK�A�
���Pm����^�,*Ǜgf���X�d�u�;j����	�F��/Ed�8Y6eYi���U^�[t�_j�cD��W�!W���2}�,�
����C�h��7���)�������
�����Il��(f�$��x�"n�������`����
�Zgd�rg����'����"�p�2ˋE�_� �J���o��Lվ.�!�E/A��vڐ(�TV�?�MI$�l��U��W��i��, �5Q�����Ff�������c��Qw������ޘ`���y���]�&8�5�����QQ!�������0{7>��P;���]��_V��BZ�c�:(��]�|��i[��&d�e�����i�@1	�]�>k)�&�?�|D�Zׄ�]O�cC�!��A.?Y��-�?#9�G��*��m&��d���RsT�x���؏u��2�����Da����%�i�~j0�5�>�`�7����	���ɲ��Am��T�Н��0Yޔ��,ӈ(��艡�L�T��+��"�]�3 7C�]^pY��V�z�͎K%��9&��݀L�ukY�-Yn�Ӊ����ya��H̿��Ovg�n�1�X5��0<�;|�J1�p�q�ϯJ�6-�����d/�P�V�(����r����dm��|���s��ly�`�b,Ͼ�5Ey��<���9�M����/�e��3�R��L�V��>���]i��oy�%;�I��!GI��tf�h�����<�	خ�n�>����1�{�_���Wǝ��{��Q��4�8��$�|���bl��,3⨞���aDbǾ�Ѫ���9X����w^6y����d(��:�aǅL��,Kuǧߵ6�M#��9��J*;���?��xw�[+�}��?a����5d�7���ৈ������Ǽg��V��#�Y��lU���@�F�)��*|��1�)>�^:�Bi�(��iK7���)� T����ۖ��� �~&:{L|���po؜����X�[�^�$Y��t�nA����4J9*/��`J��G�Ff�V�3ż�̖Xsޙc�R1
��k�XVp~[&T��b�-�um\چ�'"戤NY5�%����#�i *e�j�>����tY�F0���5�?�J���)d[�4��X'8'�6���.���9�-褺�B@����~��拵�����xV��q���/�5Jԛ�E-�}�D�?m�6�?�^;,4@�J���C�ٗ�8����� �\���L��a$?-s��ˣ}�j���� Q,�Ȅ"#-m0��kh=�f��.��['Va��7B���j���N_^۲4������C��ZBQ} �K� �l}����y��B��~P9�	
���K��wJl-@�#���V��}9�x���^eg�_����g@Nx������\����3�������ơg��8�@��on������U���R�K�S�wo�_�)�~��L�y�=d'/�g/q#\j956�=3Lg���?��pJ	�^�>-����ֳ`�.���9��npnh�N��=w #��p�]�6���&���$��#I�LpCl��4�6��T_�҇�V��ٜX��G�� 
yI�JBx�}�����R����uV��V�5�#=Gz�bC]�f{�9F�{|��	'
��� ����6 +��waq��x�!�ܜ�.�{�L����H�ҒH�jWN�m�WI)�:��e.�c&��W|;�`�2�J]X!��2�� ET�w��ќV�?����y��?��1sz�17@6���K)�)���K�\�b*�o� FU���D�+��;��2�� ��d w�Q6��Nk2ǆI��:hLc6���a��y\O��]%c2�'�)
�.|��F�>����������q��/��z�Yf	Ͳi�1�QJr���>�9"�m�>��+�0D��,͆�I�
��Ǻ�cmj+�� �?�H72��4vB<��������G{,l
Ԋ�=ǭ	£�Qˑ��I�G|���_��e?�bCU�cTݞ����#���PK��uWkD�5�\�K�wN\�Z8�<o�K��	Q�G���%���^a#N�ӞUM�X%l	���x��bX�pvq2ɫtG�̿JM/Gن��a,����ċn���I�:O�!�'l'%��I)��ᙦ��FG��T-�0����_�����$I��nj�
L�x�ʥ�.1M4�%�z<�4*(Q��d~�G�c�۱�Z,=�"����j�!�H�%lu�U���D�`%�a2} %"��gV~�k@$�y�2�����#U�{k���|���f��BR���Z(�?�	����S�����w�h�,7��Y˞�xb+O��6?��u
A�>Qh��LY��O`��_�h��aBk��wl�R��<�.O�P���,�	����Lh�����!Fs��r��XA>��	����nU~Z6��l��ţ+�G`ѭ�FZ視xF%{�JJ�#߱�3���^�������)�+��zM��P�s�������Q~:�Y<S���ÿ��C�k�x��TY��k?��������u�B,sL�򇋒�G�fL�˹���Յ٪���'\#�y�5#+0��.|d��$���=�:�=X?�#.�1vǠ���K�`��7g���B-ҜX�?���>��im$�U�Th��87�:���A�	�b�Hƴ���Pa9	��ߞH���iG7�"�l7Q��M�c���2�d>^R��[���<x�K��1��y�)�9F~v�����(�7f;��(M�Dq�cgX`�܋�1];�8���Dv��$���(��,mmnO�)߯Ώ�|VF�p�8��������up��z4D��25V#�+��{n>BdIL�˴u.�ݾN�7dVEk�Z(�%��Qb�5���,,*��%.ɵ�Syw$�tTW�H!]�]�1N�	F윅��1�K�p[�e=K�x�nQow�փ�����)1j��]L�!ZY[P��N�]޵��-�����X�VK�턏cd���#L$Vk��#�+�8P��ZH|پR!�å���V��qlZ�������qچ����6��ΨN�fgi0`1��_��g�YE�RkF�y81^Z5�//�����dDA/Z���q(=�z^f����o9��Fa͂ى���ܘ�z{=6j�?������	�	�,Kl�.��vp.���x֘Y$��<����F3��+,y+���S[��"x��N|e9�p�?���s`}�e�04�����Ve0�z»ɀ�J��6��=���u�P)�E��*��ro�.���� ��w_�c@}	������H�f
XvCr4��fsрq�]��b�0�P�j4���e���&�F���r�`����6���WKiL�`����_����ș�|���	�od�6��HD��>�B `��v���G��ނtb�F�LxÂ�$�8���8��왋�-	z�e��V΂G$�_��nϨ��?�����c�	Ω�Q��?#g
'��B/��̳�y`��TM���q&S5��5C#�U�v1)~�_^�Z�����u���#�s���� �!�5�2���,�2���o�ٜ�+ǒ�7�P�S4�sv^�h�~b�g�:�(��RZ ?��_��5a��Q�݌��N1Z�,�}7��|��s�ο������E�t���	5���e�o���~2�p� *qMSbpW���rS��{x��ftg
����f�2�}�Mnd�'���e'�zm�#�>�ou�b���P{%�#;֍-�5v���8�븗�u���ǆ�`�Ζ�q{�Xug�#��t��*�����y� %��[���!g%�̉F�<�s�:r��O W�U�(z��3�Jj
Gv>�^A��e���zǾ�m���u%�$ĪW��|`Bb'����f��yʀ�������^h^\:�i�v��^�� 4-J)9Wt2�� (�#�%�v+F�����n:Z��{�A �_�a�(Ae�D�w)�����0��$���@��KFt�؍�m<�h�p���	���o�b���Ap��q���\ֆ
.0�>D�v)�Š�ͤ�Q������+Z`���4�x��4��3�`�r��́41C���%=�h>+&�x��T�G�\�7M#W�3�LL���y���]�N1��I��-� 5�^�G�N#D�q�v��U���UVهG{} �yΨv}��� �ŵ��pW�)�]���=���2�j�+°cv�?�Ŀ��>#+;�"�2@�rhO��E��"���aMۏ�A+D:
?�H�D��.� 㮴d�ZV@$B���_z��t���]?"�7O�@F��ؙ��OFjPhZzaW!�O��1��Y�9��Xt�����D�VIb���{�V|���Ǿ�}e��a�)����p�[������GK����Q�z�_b�[�F��X�~[uwkB<V8n���/��%6+V�D�٦�}r��&�ƹ�^�6���I;xa�	��T�p��{M�x�[�٩�^}��)H=k��HB�x	!R��SUL��D)��"^��&���u5�;��g��q)��\���#�1�z���֡����!�6��Ǽ� DR��F��h�?�A�KdN�p!���CR2b�0�����f���Hi�B��G��F�$5�T/?���bg϶q���ɫuyV,�ّ�t��@��k�mADB� ��ƛ����ݎ����$�A�7��} �$z�%4�|��v�A��j���v����b�bƹ������}�H.��-��@i�So�@H>�y\/��&�xL��o�r۰F��������)C�փ���cY�*�"Fz�8��wk�T������PIFm�o������A��&F�i�1��AL������yvb��п�� :� 
˂*FVY�
=9���	\O-�A}�hؐ$'��o��	�T� ����>������qj���/��q�D��3o�G�K���/�_�8Z��M��U�nd �f���o�-Aʻ��bP�a�v^e:U��Y9�qa�|�1�L�5�{��{����D�+#�]4>Erlk=�jK����bг����*��*^��Yr�:/��"�8?Ԯ��(�=+9t�I�8V�,���Г>���O�@&q])K�%��>�n�λC�0�̢�P:Zd�����j��k���,��+9P��cc��	i?)w������\vQŕ�V�_<~�J!w��\�HQ?��3U`�������M�9s)��9CP�>�y�c�sg.YD\��3���.Z��P��_3�<@"Պ�����;h����Z��N�J�h+�I{Z8^�8�&|���Zl��W��{-���S��P����.���鳌:}��wR��QD{��X�:7kVV�W���l|�F�ۢǸ�uH�r͂���vz@�^����~LT��̀�2֑q�w���m���^���0R�w0�T}�*敤�/�"|�c���Ln�
@r2�����ל���iof���r`�%��+���Øl`@�6��|��]"�~�B��K<�94;��#��8И��z� �o�'�Z��{6����à�W]�m8��g fR�bw�͌g ����Zh������J���#��ʛ�i	c�� ��w0,���D�`�<��q�4e�ۥ��c�A����_ �HzJ	��lk�կS�,M[��d�|g�Nf(��=��I��~����VJC���B��Z7�;a�F���<���-�"V��mU��/�Yf�?��`d�S���xx�_��eW���r�Y�tJ��%�h���{BU{�kM��/��-I+a��5w�6�����*�pc��X���2�\gГ&���<L��x�ţU�9iPg1y�y����y��D���x���*A�<D�i�q�1v�~c�L�S���iu��)/`��(����'���DO3 �}�C
��h?��|��G����_�ki�,ٻ��>sXR�YLw�hI�I��xH	e����E"���֍��C���m�8��-Y�j�"��N������ǆZ���,���۾�TH0�
��$�[�q�4޻o�	0`��zƲ���/gġ���>8�[$�rAȿ�l���Z����8Ne����>QM�i�����غ�1uOE�]����l�0�ԯ�Yp�Û�����/@#��u�L������s�K&�G���G�)+D�w��(�X�s����|��_���O�5��U�'����'\����>���R4�O���z�=��?3%Di@a��;��B!b]���
P�ڶx���w��]�D�1�q��-��
=�����L�� 'ɽ�*C��!���w@e�|��Zu�,x�H ������c�w-�gM��,��ww @�U�S�rw�C��F�YT~�P;{��:�	��Ֆ���wV�w u;F�/�Ksq�����ER5C���։��rb�x�o�䬜B{���X��+~&���=o�.�^I��BD��<7�r�W�Y��Ҧ|��tmպ�˂�?��!g��je��w��v3Ͼ>���|��v�yH��o	��+Ƕ��l��\�Wwڝ�����q���+�|�!������Y=�u�?�S�O_�v6檠�����|���VV	���yd 8-��Ro��=y�]�r3C� r3v8��3 d�o�C���:���Sqk������v�I�G{/�6�C��b��EtVu�W[�Bg�a�&�U��T�{�����c����_���@S������̼	8�����Cq�}���[q��N�P�F��'����"�QD�:s�X볍\mB����I�=k!�!Ԃ�<�]óՍ<,�]�dR�9�d���nY�T�$��8	����5K�),H�r��h�lj���U'�,�>�U`>�	�za7��)J����\�r�I��;sJ?_��p{��6Y
'����67�!I4� �|�<` �����AB(U�BPA�҉w��+�S�d��w�u�	qzۻ�8HB�m���({J0�:t#�o|e�
��O�`�85�A�/�5ǁ��K�d��A�\�O���N�Ec��rd��86UP��"���h�I$���y�-��ɼ������Bo�C�X���+m澯~��[ո�0�_��AV��L���+��0��e��&�c1rſ]���\"�|I@_6�-3��c�y��J#H��b�M�t���ը|�`h��G�}i>.�\Y�D\� *2$=CBY���-��YDL�p3�\F]�H���ȗ@��CA��~�:��V�����)���b}5д�9�k���8[����> |��`��++9�1�T�Q��=��K'{^s���/"�@yr�ENn�閥��� y�g=$���wD=K�h������L�T��s�� �IV@ZL��"+�=�|;F�j�1��]�2��P����r��i��%�<G�+߼o�����#\P 1�3����#�[�0�\�!3S�(�Q��%��x��Ƴ�7�̽�_v�����2Ds3�j�*��y:�88t:0X���^�Y���u�9�o Ջ�����X4f�Y�������������WgJ�ઍ��{r�D;�O�wk9��5��`��	Mw�6�s�:���HB�ÐG��h���ꃹ�9����خԟ�=X �/�~+=D�ޕw�ۻy��nO,��7�.�~��qM)Im�G�)��?�� 	�̩��g�:��G�~l��*=.���^�	�������m-I2�aEk�V�ZjQ�SG[п(��{5��fyO��x���h.Hm�IU��NM���'r�R%L��y,�S(#7�5e��eۨ��N���Q�3�}�9a��Z{x����NǷ�Y���xZ������?˩�g>�徆���J�h#x��Y7b��g^6��ֆs/׀�[��G�~�R�J��M�	(��Ȼ��4Fn����<�!V,���9��16�GΗ�;�mK���D�2&6�i�lg��8|�B��
�A'���*ak+\6)]�&�_6`
ۂ�uz�,�}i� q�N�h�c@J7E ��:f���:|��qK%�Q��ii��D7��^}1�j��}�`{�m2*��5��M�Zg ��Oc]��q���Y+�Fcj�:�b!�R1H#��X%fU?8�f�Nq�*�v=��9x����	I��Ȑ�P	w3������V������t��s)~>ܦ��Q���ьk�l��@�@SE�4�7�/u��}�v�e_�KJ�|��'��^�_4�%�_�~�G�a�4�鮸����t��:�z��A"�_@r{y=�hM1�e� �;�_^�O7Bj��`�7k���>���ChA͎��{S8�H|���(�/ϑ��hr%��"~X��CZ�&��2���S��.q0O'��sN�ޙ��[*_aS9��v3�����[
���CG�X؁a�e�d3޶Y�g&i?A�97����(&6��h��G�k�����<IjÕ!*��� �>h��OIcNb��t��ji&�H�jz9*�%�����)���O� 	�h��1�������gE�
d�=>U��ʢ�55�{t�.~��C.roa���)�1�u|���`��@p�����D�8d1���Z�tz�S�(�@_Tل�°�'P����&!�iiZ�n��Y��gI�ס��?h��<F���jt�-8��)�'������`�5��7�Y��WābI�������9�ÞP�ֿaA�]f��.o�ȱ N�[�`�_�Y�$0a~��Je�)���֒^�M��������/��P~AC�}��"Ư�s�XI4ۆnjC@���h����t`|VeD����X��,3���:g���fױ�*Y�bt?��z�Ё�/OfH>O����w�f�-�}�H���XM�xѦ�p�60�E�e����B�T梏7Ͳ��;��2:;F���G��܃��UH�Y]SU:hn����QL��"7��2x�ŭ�W�X���*	ϠC��SDD�
3A�VD�`�x��Z�u��F��遝ǟ�슪�z��E]X��������Ȍ��8B J�qZ�x�ⱈ���r�MSe�� �,��S'��RW`��\n�N^�kg�B���5ܢiDF��ꈙC[+կ��L��
�S�:x;5̀�� ��-P,����"�g�}��f,�cR
�Bwd�$����^{��xQ#YRn���$|���fP�7�;r\�9l��݉� H�]`۾ Ϳ���ds��Z=l�����}s�k����]�~k���1��.zf�c�O���ŋR���H�)�ѵ;8Aizl�ژv�����ӆ�I�����j���?|�6q9ؔ�PEzHQJ|��d����_��Z�Q��?SS��C����7���qӚ�o��g�O���l"KZGO���gP>�pe#$Q$��]����Y��Y�P"��>J�.x���^�2�+�=�p�=�qgsU�|Y\�1x�?w�4O~+`y%���P$۴.~�ȿ4���x�}���C��,{��|t��9�hF�N�ׁ��I����8�����U	mc�������#(n�tv���ImZ����j���ҩ-�m��=���E���@+�5�����tV_������Y#�#\
����nTp2��gB��(�v��d�F�>�]�b�@w�j#�d��쫡��YV�	uN��y+�Î�_SnR;c�6��^�U��I�p�FS�f;9�_��;}��6\BP�O�L�����
_L��7{}G*{�D��c(�p��L`gbb�,<�X43"-�Ɍڗ��i�=jF����P��R� ���j�j��܅P�uan'�WSڎ���H=	,��\ʶ�Z��|,f���!IP/?T�C\@S1�[��X�Gm�d2F+���1��h��n¥Qr
9���4kTi�+�����Uy%�m�s��}�I��i��s0����4�,v]Єy�e�c.���1D�:�s<�NY�1�d+��"�D~�T��{2+�~b����O��ӛFXhƾL�#�xs-��� b��{<$@l3���wHs��֝�P��@��5`�j��9��w�f�ǜ=7]�s��FI������a��C�y�@0� �1��!�� nN��|��u��������2�)(M�����f�S�®nJ���r�%���mO�~E����ɋ��������+�~�_�N�\PQj�;����y%���y���� ���.0�v3d�?|0� ��4�͜(�,�t�z�c�z���m� ��SZO�ݫj��]Hx�L���@t��s�����;�����M6q��VWW���"���D�_���c���ۢ�x�X}yë��%���u3%9�i��G�g�Ǝ�C*'�������Chi+(8{f�n���ވ	�2��Qil
@>��X���c,���=p���;o�:��&_��$���R2�iw����~���'��ײ�w+�g1�7k�?4��OXU�]Wu����|�\�vy����[��b�C�kҰ�'\��/k>a�7��֪H �ZN
���O��(=Ϻl|���XUT �O��M�~XЍ���Q��]� ۣ��~�-cᵉ��H��O�\n���"��Cz���4{���=��h����;~��S+��(��S�:ie�ힵ����ҩ��V�K�r:?k�C!��c�����-2���|�4�`���T	/�ӘSkD����ۉ[�xg��s�l��#��x?�{ ��|��U�����TsbGbD�X��1�$���RM���DA���5g+|�N���Z���~��΍���h���O�r���X��g���г76��cb��A��X (F���W���%U���@��Z:��$R���.6n�0��i�BF-+AG��A�!�Ͷ��>��d4�o#
u�����*����JS�}��3\��AXq-_�����mn�o;���i���O���.Ť�t�AL�>+R���Ei� Z�k��`o��X����♮��(��x��R�����
��������seT(���ߕ6��d��0�,\e埤'dٗ?9,��z��3�]^Z�r�b.�_�E9�����w�����O����Y_�Y��Z	��3B���=MK�B��X20��/�;"���C��cs?>��H��U�*�)�� �+dŨ?��Hd�z3�@�FP��l� ن�2br��:���^S\�hmx�
�0��{�{o��6��,aU#�n�?No�P��x�aR֦5��y��}� ߷���C39}�>w]����?���{���M>F�Θ��l��Xȼ"3c�EC��}�z�*Z5)�ͰK��K��WU�a5H>��E���;��2�ˌH�BE���}{���8F��^�x8}a�+sv|��&����P[cL�I!��'
�g��� �t������)�X�~˵��.��e���y��0R��x	e�B8}���[$0hM���8�Xd�������t+2R}�^�+�k�GΨL����ku~���Lx6���P��I\��=�����$��~T46���Y���~1�S�٠��it���D6�@��-�Z}��%�����%P���<�h���L�*bs��}P;�kW�/��J�N��W6��G�;�r���-e�^b��x{�u3�����)@u�|(��:W	��	N��.�'�
�dT��
��8��4��x�MFy�� b���5s�[>!�:���"m)�0ô�X;�͠1C�l�>�����i�_K��-����t�Q���ع�ԏs���xl�3h����Uܤ��	K�����\Ra����h<-W�'+L�{W�}���j!w���u��Z�(�l�;#��3�,��w/`&Q`Xs�=wR`͠O8��1o���ϴ}5S{E�p��܄�,��p#�e�� al����$�Qd�C�Z?mx3u?IϢ���|���Z__���\��^�:��_�\4N�:1	~�ao�����T�3����ǲ�[n���l�����+���r�����8��K,`g��<�̳^N�6L�s7��b�{�">I�+5잒��b���������'3ꂇbT�N� ~��~�_ݗ,ZY��;68A�%����u�����HA�D�[��<�Bڳmn�)�X*n	S���686�-�HBy���z��$�hK��\RY,�[ۖ�L�df���A>3O�k��;��0��s�B��̕���1�j[�M%�ҶJ*�M�`�Ac$�Xѩ�_	�$�{�����<�̞�J�k��91vm<�� ��Q!U��jC�j���YWF1��g��^���4]VD�/�P��h{f,��ϓ�@B���zL�aE��h��H��f�>?3,��W���P�a�����y�p=ի���َ�Po�<��oFV� �tp��z�ge�:L}1π�'<����<�5F̛�c�Bw^o6D0�1O�ut��t�@1b��?TE��2������,ci�^y��E��c�����pB�r~/��l]Q8���	�����,�Yp}๝S��H�)ܛ M�U�"�H/�
^�Jr��q��5V���W��*�'R��DM
Ԋ���P|y�~	!��ۏY���*<�^^�& �b�,2RD�aI>�?u���۫���c�N��w\���p����*�>�G�[MA"NߏH�����v���>m�#��IѹA�1jQ �-i�P�hF�
�5Choс�ye�Cq䧢:5���4$���&:����=^!ˡ�|�ў46!�}o��Tұ��PZ�E��R�ju��$,{�!OF�D0ĝ�E���2˖�� �ǨM�nC�J!�|n��������}�1j���Y����n�`��W�E\�|��E��$`��[�_@�/�V�����Kܧ����{17s717uk6���	��ō�
�Z�%<e��<7M�f ���حCˆ��IQ	lY$0>�H�����v��ē��Ŕ)2~l�?��o�;܌ObY����Ꮚ��P�m�#or*�+�ش1�7�2Ex��+��ߥ%
y(���0��7���,s��M��x/'��s�����t/��ޑ�ܩ�����Hɣ��m��"K�u��ݿ�F��^c[�������V�������P�zXQ��g��/�^�Ko`3�.<�3QYh�߲h�Q��·q�o�.0(K�VKÇ��$� �gR�W���'z*��ܓ��rל�����gN���,�Þ�1���\k^�ણ�	�5�Bq�<��ML�´4�R0
m֥EV�oiT�9��%�y����D	Z�#����˂g�Z{��B�7��S%������~NӠF�|۬��¨|�$�d2J`�����,)�<ԭ��!�Z�],����,A���c�����I��z�_��Y�D�py;T�J[��V�u��J�C�V2�ٺ:c�S;.�{�Y�a���C�Ц_�(��^&�
����U��ӿ�op�i�Ey�0���ܺ���wM�2���	��0��Sj��v�C�ίM�*��s����WhS��_c�a���<��{ˀ�T/�4+W��L5�e�Ͳ��0a:(�X��1�e�<WG�B@<�AX[�w�=�����(�k�9G]�6�j8���X�@�ߔ�&�PS@4s�XG���_�%i��xZ�Ȗ��e�{
�7�9�l,���f_3�k����t�I>am������u�O6�����I5\zo��7�C͡eV�)�4��sI�#��(n��J�!,{֗G1츧J�p���z���?�2լ=�+9i�������؋F��ݑޥ~�U�>�����@�)�wD.��y��5�r��(?�����
ж�p��#)��rA��θ,�hh����$�o��nr�ץY�~�29O��E<��&�]��qx+޿�p�ф%3/����c�ե,��YeTh�GU`b�0�&��{,�ls�u���q6{^M�$&���3,_��w�1l�Ău[$B9e��,�Ξg( ��Q�P2פ��6�|�����w#���Fe�E�$���̕�>3���dYx,H�|��Շd�b���w8sw\�#���2�+6c��G�,���+'w-G�3B\O�:��3*C++t¿7Q`��+�:�K�*�����)�WA~.A"��s�:�DV0�� aw��鯣��ݫ�M�C&X���J��pb���"U�~����4J@-��G�U��E�� �Ȅ�ee ��GE�`&`L�����T���s��[,�����(�k��Ð���ü(,���&ԩ ����]_V��0��c�j��c���f� �����)x4�`*P�R'���M"3�<>Æ��zA2�nӹ�^�u��>�H
ar+�M�L"�WC��c�`mK�Vˋ�J���y�m`� wuH��k���#qM��J���",����q_L&�Q]e�D9��:��ѡ�ˑ��:8�gc#�����}s�f����i��>ܥ�^�2���Y���ۄ�D���6�+[���zp�A t�f�#�1|�3ɑ�H �?�����"$oѠL��O��,I����$t���C3g�Q�y5H2�b��" زw���(����>b�����L�\�z*�W%����C{�d�}����rP~� E�"lͰA��fC�����a������Q*\��F[W1%��	�6N�Ǌ�1P�CN���I�:�������v�FC�g�m�A��D�"���V���ֽq:�<�����ȫ&����fQ�{{YyЅ���¹�IGr�5�p�_Z���d�I��-)񄲶g#1���<�FZ�lA�i�P�'U�H�osB	��0œs8�J�:u"�� �f�K}"��h�	}M8��D(叀m�+�13o=�9�M��������.�4�q:�����h�1TY���V���:a|dʪ���P���V\h3�(���ȭM����amL���c�t}���6�N;tY�}J�(��y=�Ņ�ݱ�τMݫ�F��g�l��=D�Y����j�L-VԐf��Y�����a�m�6���	��`�%�>r� 9�X��4׊���~5>��D�r�n�\Vj�J��8�^>|�&Rb�\�a�盛5J[̊���������u���0�ׄP^������6?|���I�Xdl	��Z���[r�j@p ���d�2EB=�`��#������P�߼I)#�����Pˏ8Y��j���,����<������Phg�Ϡy3<�`p��a9���,����#��!Nn�$^�G?�G�_�ꟐR7�A&k1����n�X.�x��$���6=H�[q��D�`$I�cCa|<�[�וm��ќv� �@�2�]���Ld�N�1���<�w����+�B<��j��WA	p�&���/����%�a���*/ޗ�J%OQ�-e���XR���7�%��"�eH
mt7�j(uO�g�s�'�H��k��j�_qzɨ��?9����Œ���[�y�H)�X����t��}�5�����uv��ʃnk������t�KX��Jamu��R��1ݳe#\q�cϱ֔4��&p� �V�(Kة�a?B�M���0ڌL�dp�,�6�֮͘2�d�6L����A�>�
}�ŝR�̫|t`:N�L��o�Xn�f���4�t��������V�_��]9��U���E��aI�`��9IYC�E&u��-]U?���߹�͜�_�)�fp�c .���N��1��q�-��v2a����?�r�i���d��ߪ^��ҥ8,Qг�ks`��|E�5O������&�с}Ϫ0	��ݡK�w�vJO�9�x%�q�beQn���R���ų/M�n/t�c �s;\X��Ż�=8���r���s/WK���6�e�����V�d�̮���1c�9#)Yaf*{` ;���,;\�l���Z�5�Ф+y~��u%z#��#����^-*~�����G����'�O�����5�.�Z* Htt�Ĝ�����bt�1�2<Πj�B�IE����Ծ ^%�8V��9�1��|� �D�%Ӽ�3��ԑz8%'�%�1[Oc�
�)zw�� ,zl����"p_S�o<	�**��E��"|��b���A����$�.p�r�(�S�х�8�]�мТYU_�1���V~ =�}�pV4����+�T��� ;��&�jZx���s|\�1������ZDI,�?wCL��25�tSX��t{�=	c�2�X&V��X�ͣݽ�w���7֝!�X���U&4J���vr`Ϭ�_�=[ׁl��#�E���� ��sғ*�q��w���}T*��L�a�%�
JJ�� M�a�kч�*�o�z%�280�H�r�Ĳ����)��3���Kfsİԣ4*cIl���O]�h�#�F��@a��"���������4!�OFapƺ ��;���mf��XM"$�����W	�Tа���/���Xq���b�������A-gG���AO���c�V�ʸĺe#�0�������*�BЄ8y�ҡ�'��&�4��u��%0v��K#XH����Ez�w5�JD��>�ٚ�gs��0x�t��0�$l����cض<O��n�6�:'� 8c &R��7A�������3����]2w��ӏ��l��z�u�Ǔ�x�����Co� �F��D� ՅA<���4p���0\���|h�o{#y�J�����f����K�F�@R�C��nl}�<Z6�F�
9'��(F�L0��S^��SJ�s��FW��hH.`F�����T��s��gţ���@����L1�U��Å�����������%4�w���{ �����+A~�<_�˺�T�k������9���Fƞ.k���[ ݵ/���`��rm���5�$��(}�@{�m�߄��℘�x�6�r��h�n:�����&��yT;C3dHp��\��:{� ���
�~���}S�Xt��@�����Π9�}��W�Xǳ( �X:(\J����:.�m�gb��dE@���;��h"_�,=�!x�z���&�Rݷ��"O�U4���"���R��ɋ�Ȫ26,Nj��ߐ	`ߘ����Q�CN&A)N��õg�O}��4� �FW�q��k`6a�!��D��9q�ף_T���h18R���F���x%:����$�l� ɺ�F��T�qo�A*���/���Bo�3iOq�fT�X������$��V)*z�8P�1��P�	�K�&���MZ��Y��`L ���m�k�����f7{&0��~�u�@�[��G%������˙G-5K����^���q]�2���^�1�(PE2���U.��u��g�00��=�s*��Ix�������$�y�0b�>���%,��ËE~g+��{�]����<
癎����h�V���1s��|ԋю6�+�5��w�A+*�y����
�:�_��D�ѓ�;d"�_�^ft[F�r�g��"��}iOhu:L� xf�d`�0H��A4ҝ*1P�\'b�4��Ցb�&AVn�`�����2Ⱥo�@	�/��8)��t͂�%�vC���lUԪRۈ����>���x�X[	�w��b��aW[&���t�nf��]�L�}PS6��T�&S�$3L<O�)��V�c���5�7��*_"��БyqWb�F��	|�h��M��d@3���<�f@�!҄���#�k}��TX5Y��������c�ݗ<p�����/��>nAco���'�з�"��GK��h{�cо�u����I3�� 4%I���	�9t�խ��w�cx&�����|�]�]��U!wb���C��p��(��w9X�ұk���l���%�a��N`��Z?_�r��*��+�1"�fh��>"����� e.��_�u��N$&�|f�B�����W�	�Ҏ�*������SZU~Ierz��>��C��Y^\��?)��6�T������E��f�"j|�%q���t���W��@���?���d&
!XW�lS���e����,W��b=���d"������'�
���,��!JF��}6�gl���?�	��c db��q��Dǈ"m�K���~�q�C���J����W��)�U�-pKH�胗�pQ P�͙2k��V�v����$cT��x�/�rq�f_�B�,g�t�ɱ ���.�jmK:�R�a�^3Mc��-�V��|5 ��KX	�Q�l�ȝ��zk���K���Xx̵�0���!� �b�ǁS8�
��#/$mSIP'�en���&���nX�	kn�i'J��/���ٷ�Ꮉc�NO�vYC�!C$;nk7�b�z3q�Ĉz�lw�,{&�k�g���t![�/8l�#�f�FO<՞�b1�
����K��3�����
N��װ9�,�8�*��lbK�}�F�t^_�s���%��p���h8��1�c�#���@+:��)�ҟp0�Yrh��)U[3<��a7�}��%�,��؈���n�&��4�B�}�M�*�|��6V<;-��d7GB�u���&���/�+��Ha��#߉�^�K���(�!Ӊ��5k ���b爆ϡG7'�aWV�{�Y��#�B	C��;<��5g�g��/��u2J&��T���@���E�[R�&��/�%�{�q׺����_�ӣ�y�%`P�O��2����0�0^tf ��ܶ�؅�a N�����Ƨ��٧����!L_ׯ�\OB���0����Ɨ��iX�V��G�囔�Y=~�QQq����3yi�&�F0n�#���*|a�8�]y���Z%���NI�{��>�D�l���@�)�ԣ�[��d�r�-Z��6���3v`8��Q>r�SG�l�aK�(�0��)Үd��w����(pgʿ�B�0���-&Ԕ껳���e�&��b_hęm4'��D.��{+������1䴵@ۉp���c�&׳�+�\��?�1���|��u����`7]���XG��2!d9���F��}�����.���Ώ.�/@�5�Ձ����*�����5�R�M�qiw��� ����(�Y���+�9�i3u���Rt�'��5�B�nOB���Bt��3b�Z!1��ؚ��s-�7�Z�g�o�PS �ĪG��wW�m���]mUɐ<�:�=T�Tr�����g݀�׿��հo��=A5#��ney,F��#P��t`��
S����E'�H��5�ᬌ������?�6J�{�~C(*<�/_h����\Z-L���!��~���0��6�q`Q���g��i;:6�D�\�<@�ֿ�5����_4���/4 -}��FW����b��=;q'6}9;���!D>����V�qLr*ֵ�ߒ�u5ၺ�ᝥ}9����4�\�@�[��xd�b�ܱ�Z�:-|��:��eA��_�"<������`��q��_uw=~S�Oy���+m��w�*�A����ڳ����A0�&K]�.n���ڥ���rt��tZM/�&���4�����j)��pn`�>0��F	M�!EA�1�c<oXű�S��}Qm�K���R�:#Ȧ��4����'�2Y��A���Z�q+9�t�k����<E�nfB�%�)�<��G�=$%�ҽ&�f$�$g�a_Ŭ���F/$�+ C�ƿ���U]�'����9e����m�.���O�W�{��3t~7��$�C\d+�����%6��91��>���Ub��&��#Ll�k]��tS%r���C�d^���B�D���/h�1Ϯ�q9L���?HX��۬C���.�H�v����_�s�3� �X��O�T��Py�ӷ�/v�¼v���;��a"ŒT���ԒE����p�wG$�%`�Dt���w����zČ����m,i\P�X��=% �)�hX�m�Z`�L9����9W��ХN]O0�r� fS1��<�ކ���
:�L��ձ�L��1&���ߌٕAH��!^��R��n���(��F�(\R��vY�r�E��Z��R8�a�}1�w��Qn�o�@�>�NT��49�S�c����I~. �'7��4�)��S��wE)������I��"f O�XQ'�ۼ�5t	��Sk}���;d�mHO�6��za�?�q�d9ݰ�+d<�(��Q�|��Z�C�n!E��}T�뻧ٍ?���zw�AJ�����l7��?�zG]��98Dυ<��}uˠ�|�d
"0�=�VZ��3�boF���M���Ѹ�:T\�
�-��t<��QՕ��8㱑�,c�R� wij�}����ڐђ[AP �*�}k��͝F����v��Ia�;_�b���8		Z|����ښf�EJ�O�/E�����܃z�dM\�'�k����aKi��\˩�$q���X��F�^�m�\ȀthN24����H�7�7��&�8������҂�K��"�=�*O��hQGL����a�6=}�s��g]��,��,���P�c0�kl���k@�&^����ڙd�T�`kh���lp��� K�����
����	���*	RrZ�y���-jkDq�Ȳ7�;��͏����
/I_x��C���A�g�zs�xM#O�@���>.)ē�ˡ���}�.�P���E)�G*�����8�H��\���cmi�2�`�@;H88���� �gw�-"������M[��Լ�r���U���ޓ���֤��>�a�a8%�_�J�b�˅�C�������3/�a4��(e�X����"wu�gއ�Y	#Y�����{���KhP>!�
֞d5!N��`��w��_�W��CWc�7����X�S�Dq��Y��	?��� �B��w��q���c�\+�?}�ۂ"t ?��<v���4Mak8�傠�0YzV��i����e�q�I:�r�Gb5Ƕhce�֕�9/�:a��#��w-R'h��k��
�έ�^��Ƽ�@n��b@��}k1�
 Z}��ʾ�3�a������
�;��H��v`2
�%����G�%i)���4���_XG���qn����/ ��=�`��B��'٫���pF�_�Ac��w��P�}�f^�?Rj�~=>O�3yJk1|�֒x����O�8��L�f"��\�ƌ.]Z�&��%s�A������,�Y�e`�_���)���=��yeE�~��/���~
&�O��XD��cF7������d	~*���	�"���-\6X���h���}������۠{{�+��tMZ�F��h���j�����9�J��5�L���2A�q���|�w�6��Ï>�t�?� xIT�xZ>�ԕ>��!�O��=�:�G$7ɇ�rؐW��"��{�e^V����F��Ha�a ����S̴#���u MV����^��,�JLq�,WM�-�{U,ԇgw������4פ�nǎso�R�9��(�Ք�h�?_��q��]Če�:��&���J���5^To�<��Xm�/�%�Α#�Y%�M�� a�,�2Y(0 8?�;[����=kze�S;��4��a`UHu�\�V���60�M�+�$Օ�',
�"|)����B�c!��L����L�R�ʍ�""�T;�ɬR+�	߲��ǝ���Hsy��h�-Зbl��-6�ڒ�;�� ����q �h63@�&�z��;UN#(ht5���o����g�8a��gͲRV�L��"zR�Q}la�S���Â�G���FV�:���|�p�gt����0�U	��)�x)�c�/Be�֧�na,�FS��������T�"�a�r>y��؋W���	��m��v�.��y���Ao�J�u��`,�ۊU|�D�+�6�/��b�>M��i7֘j mVY���(��p��/�C/�R[�W�� �'aqC��{ 	�[&�5��� ���i��ˇİ���D��8? w���q��`�:�����ܶ���=�f��"ɽ� a�fw��Z��uƲ��Z<E{5��Vп�L"�$�$����}�D����'��)���h�!N@�'�s=�bh��n2�����'��i�/XIh�!o���y������Ѡ�[�ﹺ�x�����s�NC��~bM�0�H�ay��@0��q�ѧwm��]�G�/��ͭ�&]�� Y���%�d�0x?����z�M�e���d>� OD�D{"�tUR���)YJ�Ϲ��d	�Ĵ��땶&��H>�EL��q�������H*<(�*T�6���dg��/� �l��6w�;���A14�xʶ[
'����4zQ�+-0>�27ұP����X��p�|h>��)�R);
g����m�a�S�\�<a\i�n5SV��)'G��D΄<G<�o~HQHjCs��>22���Ow�i��z�n=�����L���Fl�X�G�d��F[�JnjgQ�fn&9uj`dpıH�7�-�O�rH���>ܼ"9�
�4���qh�'�q���v�rP+���y>MH�����	����t�Z���㍰kfE�lj�(X��D�}��J<�Z�Z]�2��4� �L��'�����(���&��M1�%Wq!TYg+�˜A� ��g��,����L��Eا������"^�,��({���h�;Jj����nk��6���t��!v���Oy}�&�h�?-�)qY��w��}��.�O��/�Ɋ�{(�K�^=~|̃�����wL��~�%��Q�U��=CKΧ�id`0�]Τ��9���I��_�gL:n ���� �w�9?٘!�����	�x��I���Q�J7�>&C.��ڻ*��Fė���D��'�pa��8��hl�O>��qZ髈��]NW��� I���>+a�{L�0���Z����b���_ީ:S��%֐,���bT1�@2�69]9���[������� �����Ԟ`sg9�1�x����;>�H-�w#�8���K�Ĵ )Ʊ�̥�@뉐s�V�J�z��q8���z�o�|Lz�;�<����)u��g/�%�}ᾙ�N}��D���M�� ��Z;4C}�9��1vD��- ��ߒ����`�^�H�6;�s� �`����Qk�RTh/�߇�Vj�&�n��%ɶ��B�c/"���FI�4�eZ�
o�a�H���{���q]%9Q�b�u��t���
��9a�'Չ?�ǲ��O>0@��]sN-(=�[v�����aB�Τa�T؆b����)�>�sU*���0��&��7 ��hk[���Lk��-T�Y�+7����P,zSV��X�A8��ɸ�2�\W1�z
 ,�ؠ4�5¥��S2������X�*�G+[%�!�_�$��"�\�5M���W\	�Z�*\�����hF���a�gM=I��g#�_��5��sC-���E}:U��L*��VW�/��H+�td�W��	�k��״	�U��gJ��~����.��Ꟍ�5����_n���p�=�70�wH��xM�#����LA>�E�s�����&�n\<�h-�a��̊���Q���L���o|h����Ә�$�I�vu�Hn�M�5�����X����C�(�,�P6��uL��ʔJ;���*���'[����W�)F5����bl3	�|�g�ʻ�����bM��]��nm�=�,�*���n�C�#��Y"��>���Q������-�T���b�*�a���]��D�Lsռ����[�[2�s���&���`Ij�Ow򳹭���E5zR���bE=��#m�	
�x�ʭ�2i�q~_�Wˠ9�%��!2%Etи�xLH�D�v�7����R���H��K���ڶ��W���FG:7).�ώ��꧶;��o��A��O����n6�I	Аa<�b��y��� ��.H��=��t*�g
b����D�}y� iJ&ޱ0�H��Nk�2��R��f��EԌ�#ֲ�p��}��k(���W��^�c^����ls��|s��ȱ�y��ݥAJ�v��C4��A��cP׋O+�w����i������2n�O�nJ9I���W0�K?�%��{u5��tj'��*�d�]��̭�s�_l�EgW�4�.4n�	�`�j��J�O�9���Y�[R..?���|�޹��܅�x ����<�{��v�b�|�F���(&u�`�\f�~Ɛ%&-�`$|����5"�(Gr���RD̫���&��
��QfƂ����� ƻ�§��z�(�X�C�_�!+�,Ę��=�;�/?��h�4;o�'gK�Ff� ���=$�s��� p�R�W��dвߋ��jZ�R1�I�
�ySC b�j&�+-�UP�5: O���yw|Ş�;$nO�X�uC^y;�vK���~�K~��b�!�羛	J1K�	.A��d썬�R�)d<�b�$�H��^�����PY	�髳��;R׹�Ah$n��0����l�p$�R�Nr��`Ի�"˝��	��O_�0�>�&�� �%t�
G����8��X�čE�{{�	\�.�P�4R�t|�a�rl����� �I��J7�*,��uL9��P���r���Z>�E�an�>�NeL��J�����Ĩ��!�}7I��e��ȳE|I[�2���*�BEp*;fW3j�}�����<������^�Ǜ�	Wr�J�`�2�aAިo<\�ܻ$�N��/kn��Z�Tckv�`~rި`�.�΂��Zon�t�Y]��s� ���G�J�ma���\�t�X����m~��CB�W���7�ع�ҍ��I�FK"ԫ�ܓ@S�C�dkc�*x1�ꄕ����E��׈5k��t�:}�c�}W�xQ/�����2���]E��r�s[jh���U4�����VaZ����h�z������?:q*�Q$�|�X�3,ty�Q��x��~��$�{7�N��*����`�Z��.�W�u�h$S�IeK���)�B�ΰu �d6"Ia';�w����)p H�;8���i�)Qv����[�8�穖�M�)�l����ZI�V��o��}�?�<�	�n�
X���n�4?�4K:9r��zsr5[כ}3�C�-:���1��btk��L�άj���M�(|k^����C'�lm+�6�x���=Nh�2��1�GS�q��$K�X��� �Q$;��)�����7 1G�6%����j���?Ex�i�������^���	�ZL W�p���#�u�����Ն���l�̜� ����26�=�UhK$T��g�L%7����^�yc�lF1\��Tx3Z�Z8O 1Hs�fWQ�@a�D�����9j�J�O����c���M�y��@Q��1�"�3 D��(����>�BO�e���#��$lf���	]j=�����o��Gt/��K�(w�q;P���ͼ���$��rǼ)��H�@&V��j�ڜ^�JW�4��~�e�ӝ��(�$9?;l����A>�5��j<qEA7W{�Mhp�/U��Ʉ��b�r4�(��ܒ�r�W��0)A]&9�0�� Ԕh�"��byES�P�i�>9h�HI���b�pF��f�%���d ��^=�8k��>H_�\3XDaZ��~u ��鳯����K��w��~̜�qE3J�Suw�Ш�%���qz��[_���5oB�$�����j?��3�"d�F��rQ��=m���,�@&���O���`[+�O����3�fƻ�bM<���%�U�ٝ�~+�k�i��Ԧ@xF� ���.���g����,fQv���Dڏx��hi2TҮ���2�Az� �W��&}R�E_d�Wd�b�_=���Mi����T#G���O K�o�o!�)*��[_JU`����j�_�c�i���TGU$�1��U�t����;,��³0:��v��89�SY�;�2�� �� �jGrZ`^�+�{L�`T4�-�׎h8p>�.�q��!�n��Sx�[�����ߣ(bشe������DR�@�Eg+SE�c1��Z�O��G�m���%Om��RO�iW�X)"�͈��(��ƼN��kkE7������&��X���"ʯHр�C�X��q��i�Є3H��F�2D�"�oXI
��^ ��o.�f�[h��k<c�Iφ��n�/w�rK�lz����	�J,
C-5K��G�Bk�.��b���=wvP��c1�
�h��if;�=��'�L�q5qշ�
�g��Nf�+�n�ח*o�լ�p-��<�˫� ��`MXE��&�TP�B��0��!��8��Z$��@Hk�����-�s~x�(Bp�Q?�5��iKee^��D=�}[N#���q,�;��W��0L7�A�QC� !j����B�t0rw�(�]Q�6!i�7������1KA���/͵����3&�k�������_���w�3]�^�$w ����`S��/\%�lC���b�V��*2WX����IrT���v%���|G��U�C{׿��uoѵ�"��֠�8�q�K�����G�s��HWJ	��u~k�5	=�@N���r���I�=dKlM��Y�qD�غ`�	�W�S��+E$��7�!�ʛ�Hy$���*K��	3�\:�>��$�)�����s�L��6';�?k�<�����\�V�1�E��5}���〱�B\g��7��P)i�\Z�J��Ag�d��,�w���������}1#)8�/d$:%p1�G<^�S)�	~�<=�uJ[t5-�F�lQ;+~Q��;�_��A��t��aH����G�B��m�D�{,n��\Y�3�,���@�N�/]$�]�*�dSS�;~�>yG�z���}�p�t*C6��~?_"���6Nx���tj��i/�-����V�ûNݙ�0�A,��,@�0��,\j|!�M�P�Oµ��9= ��=��x�t͖-��L~[#����Qls��l_�kJDp}�4y�k��y0H�����$!��Ta�2��0?c�Q��%�[0�*�n3hy�Yx�ܑҩ��2y����{�~�݇ S��$��N�?��#]��ޛ���o1�5�{Aq[7yA��#��[BrO��]�nk�M˛O��!�j�@	9?s���F���#d}Ml��4ؔ�W!�z��[���q�b9��W�lU]΄�$�ƅ:>��S>���NM��B���AmČ[Oа	G���o��<2��V�!`vY@^�ϰ2���z&��!'>͊B�U�hP�G�8h�w%f���&���Tv�����)�"�&�=�a
�1��YJ�[5�e�BV�6$�/�������	���>�� ǡ�o��*"��h���O�wk�>�EA�,��E�"t֬bt���W��)�*Ï�_��5o�×M�X�q��"rEW�/��64!O؂9�li;HS<��١���<)_ir����DO�Fg�oC�;��Ê��Tp��߳�}bl�C�h��E�Ӛ�J;�8�����Z�L�#y���܁�S5��jx}��&穁�1��Cf��{y>3|�!Y>��{^�f�������ܛ3��� V�8�%f���DU �;%�llxJ�N4}m�[Dg���T�v_IHս)�%����C����,a֡Ľ� ���gT��Y�k
e�.���~����!K��7�|�V�Ɏy�o��H�W�^Ě�t����A�G�5fh�̞߽�XO�i��Ut0AV;/���
g1�7�t��mӠ-0h<&�T�M��%��v�}`����?
�n�L܎�<K1>u�Ӓ�֝��F�[��Ȥf�P9�+ �f�fn)����2�����ū<���+ϒj��Q��Mx����;�s��%x@̼� ��2f�� ��m�2���#∋]�Y^���xk�/���8��'����B+i�)�t���Ěft�wi��-���#7���T��ka@�Ѫ�Nx�d�JoV�������g���Z��	/��c�����'�~�p�8�tbC%Է��[3��i���tɷp�u�~V+�!�����CTL}�$����M.;�}�E�#�S3���I�ʅ�Ѷp�p��),����b(��(m8e���l����\��AD�����'��-��&����e'HԜn� ��w3�7ӁHӃ��L�����ͣ���K9��-k��ED��hۯ�Fb���vU_�aF�޵�<�+$��n]����q�DW��4�(\��	!�\��j�z/,G[(��~P�K4��Mh���q�NYi���Q����.��XY����	�����J@@�ݐ!����Π�	�<�/��ۃ��mdF�F��� Ӂ,���,0Evd4,� ]�`�_��&m����*o,�y1 �̛l���=��.�ag���|بZi�lw5���%���P�i?AѼ��S���'ۙ��X�'v�^\���u*�}���t������v�I�!3�
m���.���|������n���H+�(�al��0�j�(��
�A`��2��t�p8�A� ��r���Vl*c�^��j�mu�a�L�Oٕ)Oxi��q�z�.�K�(3E-k�v��n�Īa��*Ľ�k]U� ܒ��#2���|c��f���.�2�ivSD?_�"\<3o�(u��k�������R�hW&n�hJ)�wym@�?��C/��t/��$V�V�9��X�T��)4 һ����ע�דK$3�i������yx�PE%��<����=���	���xEI���M�ѩ��-N̡�l�u���ⱨ┷��}?,�y�]E�T(�？7���s=����$�1�ɿ����f�j�~�2'��U�;A�Έ�FdS���N1� ZX��H���<d��:�R�"��.�uArq +"�&��+֞��u.PY�|�k�n�ksͯ���]��\����	��ԑ�v������N9�A��;/C�q���`��,h����}�˹�p7�.4׸3���y���d�>�p�?�����ňs���?�;��a�����:��](����Au��-H k%[@c����޿o���b�ۨ��k2jԾ~�g$.�a��%�e!����h���?Z�眑�[o\z�F�D8�Y1�bD<����W�'- A2�99��Z�0Ko�WЦG�%�䩬ǣwG��X� ���A&�3!�0dB��ud���ӱ7�2]�;B���}�����������
�(V���_����ܭ����~sY��j�U���!q��n��t �g}��U�I����j�s٣��$���,�!	VC�39���Cg3�y�jT+��9N��v��z�(�aYE����y�.cR Ё��0�`�Ƿ�<�:ʟU����}�s�7t4A"�)}F4G�U�7� +��\É���YIHq
cu��#^� gڹ\�ς0�8:�j:{z  ���-�YD��T�Z6:uu$Yp��Yn��-��FПL�Aڝ��� 
C�4�k�	vsH�?Aˇ����ӨS�>�:�9��'��/Vh���m��wh!���7I��g_����1BQ;��$�3� M�`�-'a�sro�m,>[7��ۖA@�"!��{�.�����r
�񘎢��%b�ͳMNaّ�ھ\��咬�]�U��8 ��=��@�doG�S]Y��*��%�
��ǉ%�
��}��ߕ�qyҖTJ_��|��6�j�)�F��_��ĴZ�և�� � M�~��!Hrۿ��'��P�~=E��!D�fhy��m��a-�.l��`��g�ڗL����{ǃ_7*�|�C�}�t�����@��DraU�U���n@S�ę�q�öPp��,�D���� ��4U���E�$A;��[�(ޟ0���'Xp�����:C��Kl�>�jg�Y�kR�/�
��GIy�AR둳_ڢ��1��Z��I۹�O�" F1�b.����B!G�Z�V���׬����<�<���w��?@��"�N��h�Q��\��� u�.Fu0�21l3�`�i���ֈd�k�x��>�?�-�T��D`	�l�t�Q:7H�j��>[�N�BU�aT���xE�UT� �$�˲̓L|$M$�	��+�Tg�<��<ngQ�>�ۇ�!t�:�N�1_g�'�
��J<�!p�Qx��q\x@��������V>Q�ߋN*%ff��&Лp��.{�^4 c�� %�"�6�r�0{<4U}��:�i-��.�/�P��#o�5�á19:��,�Q�ct.%���di$�@F�X��5 ����X��76�$��A=�{+pi	>�R�ԥ��MR�&c�&:���n�c�ע����NC���s5 �J _ٸ�*f�#C_b�v���D�:��N� �>��,�w[Auo"(�S":*�)d�|7P�������59q�6�:�'�L�+@SEB�s(��$��KNY�	��R���\�� [8?h�3v��`����Qi5P�U�ms�ݷt�ማ4U��]�c�� ��;���(�PK& g�*K�HB�Kg��:�W�x�r���=Y�X����7�s�,��`A��(�ߤr�1P��H����rau�Tkbk�.KS�w�6�o����ǿ�.����6����������ӡрĐt��Jv�_��sH��iC��U�:�h�:V�\x������v�܉����ML�'Px�G����,�cg��\�S윪��I ʡ��tgI5K���)���@��� R���8|���A_8��$y���Tz냘��V�~�Y�+�����9�3�TK�J�_3�Z(Ҕ4"�Ur.o�ۼBy�͢�]��D�U<���I��<۽�|\3U���-T��%mGM�q��������%.�AO��Cѳ�\��R2K����}�fh�&%D0��:�dNlOD�q��:��_�\1�]
�/��V���w���${h=�!`���;���%p��1d�2����C[H�^͚�	ЯI5�+��!-Sz��/WS�V��^J)�Z����*޴��vxs�`�_\J�f��)c:1����	�*�t�;X�>`��"P��3S	+�
t|鈈�ƤU5O��fF5�^�m��y���� dh}�򿫅α�����SSY�)Hr�4����~�d��=lᮊ]Q#�5*�j%P��ǎgz�b ���>�tr؂a��k�K���ӟP��ZI߬�%r����C��>��S�b¨
Q�6yJWɈ����n)s"�� j�ɉ#�وtS &��6&���ϛ�Pz����E�
�����A4	�/E�n��_%�Wr�7��%xb���d,���4���BM�ϿP����:ʧÆ��"7��7d�Ǵ��?��l"@A k^�B-P�ʧ?�DK�JVU�R�;�X婄d.�3�|>�e\����:�6�o�T��A��'���L����{�����աwZ�;���V����!8�e�E�"{�m^����!�]��N�"�9# ΐ?]�`��J��(���N��aF��ӝo
.��R�˼�����jZ�����#*�0'�A]�n4�b�8I\̍]Q{��B\Y��>��$�����e��y2�w��3'�@���M�0�01]b����c7��K��:���I�-��&��(�C�m��k�K�1�IzRt����d��q�f���|ɫ+�DL�7�G�x��q��n��!����[��R�k���6| �O���T�װ�����K���� Ǐ-��I{�>x����z�'!2�v	 �佞�#���Y䭻̚u'���d�O����%�S�����6-͌�N�EjkD9�������(�B�����M1��7�:��셳F����>��?�;�D*0\6v�1~�W�����A��:�2Ņ��eiL��u��*�|Ij�HW#�hqd[Z0_��o΂�gU�倘R�m�2�2�����ʛL��L֪g&d^x/E$�m5���pb�	�S�h�N��ڲw��I��oE/�=�*x<�F�4m⒏����`T#y��q�Qu�8n����;5�94n��p���~n�ˤ�4��'�Yw	��=�^���Y+�k���GJ������/��o�ȭYc�k�� ���%o�9�U�Y���ǅ���K�&F2f5^+X~��_J��e ��)X<>�E%�������K/������^|EQ���!o^�к[l��M_�"֑p(񣅨ls�\��Vh�*��g���10��BCi��Ӻ�Q<�� ���ɠ���*�������.)��$�cu�������b���UVA
Hm�3�4��a��s�3΂-��|W���L���'U����c��P���ils`�D.��S*����oQ�4���{�X����X�[�A30��J=j��<�)_9-P5�&}�I�'rXDl4y���V�Sm5'��ѻ���g
�D�KO���?Z��o(:akR�������L�|r��\��;�q�����xL$�ի�N[�4px�i��L�sжMN�g�����>��,c��E6J��;�z+*A���q��#,�4/�����[u&�_U}GnBy�� k����p@IWǍ�O`g@�_�mh����_ݼ
`r�	֑W�P72���m�D��n5I���@��N'QZ<��)�E��=v�iQ��(�U����pY�u�U������	#�`H:���U��g�D���&��������j�/�Y��Z�4���o���V@��M��ʠ;���T���� 7;0�]��Q����E�Ĵx�G�ĳإ̿�1W<�9�F����BE�r�-j��������1/)�÷6;9���ϝ�� t����վ3���C���ꨵ��)���
�t�#Y�ġc��{D=�G&�U_D{Y����j��r�B�le���cXxX��F\�e�����+kٕ�"
�ڝ�%0KN�G*�eo��%�e�-T@���p��>���V��_�k����#�߿i���+�h;�^%��GJ�j�����ZN�i�\MF��c�&�#�m�(i�Ha`����㶫�N�� ��d1Q_�60�\yA�b�Y#�x;�
g�ݧ�z�F[^�������T���
�Q6C���*��~J"<J
�a��P��MR��<��2+��*$\��p�0h�b�&��-I+8E��))�Q[O�X��o�|[迒��V]uQΏ�������Kev��y�����
K�`n���=L��ū#�V��-z�ц�蜝�s��>�$5d6�5�h39�S���c&ԇ�*S�f0Ń���]��ᔥ[ ��a�й��x۽vr��A�Ҍ�G�����0��W?́���	l{#�I&4��x�3�G�������7��9�fT�*,F�I�`�U�b_��pg�?g���{k�V3��!���yPp�v�Ӵ%��4㯳5��ީ��Ҵ&���(�m�/Ѷ=y c,�/?!Ϝ5���R���ZOF�/d&bk�-��{� W�X=:%+��\ν`#�\m�K��!9�[9�����<;q���SC�
pk[㘂� 3Ԗ ���U�SӇ]'�	v�5�ۂ�]�"-�����o�ѿ�L#):��!�_:0�0���:Pf����lݣAE-�:K�.��y	#��^�e�����X�^-53i���6�f�kv�
aُvmR�z�X"y-��bz��E�I�IӅ~��$�iRE�Dm��M���!�qn���=ټN=�`�z��:�V��M�7�ɮ�gs�HS��ʮ%�/:��	O�������X���)d[��vC�b1�	��tFdxeo������E��uX����8�7�i�/��2����MX���B�SXEEm���<�#Z�g���/��Q��>��s��<�R;����z}�3�J���BH�Х�֛��:��,�con%���>O�q���<�S�Kk�	�~�����]�Ο�_����W����&YaY~�_&}��}�ٍ�e�GU��D
������J9@��Z�c����.��;�R��t�����+��Z��M��o�Z��A`� UW ���ӹ�`�:��q:�� QD�g�-C��yj ��9�J�L�;?���}��ᬻ�HA�v1��I8�\2֪*lA��@��E	�P�R8=�6#-�ز�����ŭ5>_Q�	�E�πYF'�X!Z����j�3^�]F�7���/��X!���*��M��;����L.�	2���z�m犎�I�����1�hǷ��h:�擧���y���_��2ɋ�8xs�.�>ð���~N��S̵�)�p��+��?U�t�į%�g\l��d�X��a�%�~�����J�N��V����d�fޟ�`}0ƃ�j�z(��:P�z		�q��3�+ˑ��ť�C���&"1"�]����t��$�ZF�6q`D��+�� O��N��d���q`sU�*y
���ޘ�j����s��3$�C��2��V�=�y�ZR[���/�ɧ�咢���`nK��M��#w����tT������+'�t��|��-s"�_�F�L(Hp����T��on'{jy��񃕏R��>���O&]���q�b�_`L�&�ޑ�ң��/��n��7��7H��Z ڌo|ͷ�t$Y����ތi$�ze��-Q�mlg��t��]ل��3��-�u�Vӓg���ꮎ�$4�����Ne�׉��v�=��-�;]�@�a��ʂ��������zr��+)����i�����)��C{�k�4��ٌ�D�������FP����wu��w�n������cڎ?t�ҵ�J�n:CUi$�/_]�r�k��&��bW��Jo�xQ)T�ekv��'1@w�F*:�j����%��w�����Op˧�r/���� 3&������k�}- H�:�%G:�{��t�g|���!D��DO�	��^���0&��|�%��Er���K�a�)�e<�.PT���! 0��Io�I��۸Y	��H���, �Q�H���r�K=���9ު�v{8�ꢤ��R�>��3�Z�&��S��+&mn��H%S"��ؖ<�^H���jx?�`��`%�(�{Q�f;����u����Ny�,�#dl�n��.7�Y�r��vrU�U��&�0ɠT�J�w�xs��k_y1ܡ�����;>��ZCG�(k(�i�FHo�*`�cꘌ��]���2p�y�$"�����U|M�(� �99�W<S��f����c_������ �Cᬥ�l�S��x���S��������~��� ��5f���(��}?O,���ʽ>�>���Ї������~s���ϻ�B����`��=�'�k��b{�;Uh�������h%"33cD���?B���q�ݧ%�b�Ҿ����7T%cٰ���X����1���l��^���pH�S����O�Li�g���W�!:�uؑ���oh�g��p~W��]���,��$e�^�\�*�NŽ��H�\��^:k�L[$�fѯxT[c��[	��(�r�@^�P����(I�7�H�+�%��'H�t���zau���y�Cx��A�a+	_R��yc�s�˛�j��؂�{��'���~�xYz;!En]Y��y��:ߒ�������@�d�G�	2]:�<O�y5}3�E�BI_�m;�Ǻ6��X�b-�򂷝�����RG��*����L&��������3���K0d��P�G��!#��#Q��ZN��,��5���^��(�u�CΝ�l7g�4Wkq�)��-�T���!� �#�!2oۻ4�Jv�ɪ�N�ķ!Uxd��(��W��{��Ɋʀ�\�ڧ 5G-B�O`2(\�L�m®�|Q��Xy��H\?�&���{Y����]���b���h.��O��S�O���@�����\�Ms������j��O�#zj��!�HP�������Rkf'��	j���`O4	�R-�f����ԾF�:�<)ZXFۋ��8��N5�\�ƈ��v�"��]~U�,�_��0r�DG�����+Y�._+��E��=0�(Ĵ�x�l��+��i�˕�.Ϭ=�r��LA�+����Y��M��:`�%�_��M��dhTi��E>xܭ�JR�>�wv�#^j��ܖ�nm5,���J�?JMH2۱t���?�V\�GyiC��WWYX���T8��0^���p�c]�?4A���ǭ��7Q�D���G6����A��z���&/%zf�������bk�G`Ƅ���/��[��ooU�y�g���j��Uyd�C��#���^]�"�.���_�RF�� Յ�{	�%=_̹4n�:��ӒZA���w�vdN���B�@�x�'?���k��J~�7�"@
���#yDr���iDK�@���O��_�L	�"4����b��x$���N`P&�}�Ι=w6w��Ɨ�(���pA�6����b��I��O��
!���J4 ��QY,#�Q���`A\����5
�3��ˣE�Ӗ�m ���R�=��v��T(ّV�A*��B1(�;��Yͅ�۳.e�S��ث�+Ԅ����˻2hf�QSx��$�G�v".�����ȼ#n��z�&G�d��	p+m֮,�A<!���Z��T�H
Tʠ��6�_1,���cU^\8Bx� ��1����S���*ݾ_�r���7ˏ���g<~coxH����a�d�\l�U�� �yN�E\R����c{g�U�o�坃[�o�pX$$Z�mٶJ�y��%���Εj��_��å��7�k���-��NO9��u�:�p�N�$�>�X�1\�z0@e��%�����Ly����!�7>&�SД�j�W>�%������'�&z�ְ�+��휼�
���Ӻ���;��b�V!���4��������6D;��J�B�
����G�"���^���O���O������I�tEXg������%�ۑə���o�J��UW�b����&�R������It�ѰEv�Y<��&K�J��B!S�l
�Pq�y�iG���%I�B�O��)�y�3�BY�@C�5	M�d��H�I������m&�LV����s� �K9�ctl��,�����y]4ARĘ�֙�>���7S��f0�ZM;`��29�a���l^O������ü��qȊ���#;j*S�R�q���g�Sy!�j*J)��q�Ol��5Do���t���HC�� 1i�N�����:'�Qn���ڠ�3�8z0F����&A�2\]��d��.]��"HAS�C�|�%�OAq�8��36�X���y�$>F.�&;1B{�un8��������-�7�Z
�c� yJ��#�4�;וX�.鴦d�èn�C`c��-�q~
q`���XǨGY2Q'�������.v��id�!L=k��M6}�e=�ϥP���t>�)T7�NƊf:�h���1�)�M>x�D�v;��,��G&;V|g�AzH[ф杓1�ۅkm�w4Ǎ�B[Ce�\@����W�U���L��Dj�;d�u�HS#ۮ� �#L.$��<Q��X�|�M���Dw\v�VU���S_Wۢt�ܠj��_L!����.g���z.���(�K�8Ҋ�H�,7��u�iwKg�<�	��'�R
/ �n]�i�#ǹ�̋r�����Q�
k����2��B����	G=����8��AR��J�~a�����\ז[*�I&$���|�".��/���g���@jFI�3�x��k�%OgdÂ�ƥ |}��cޓٸ���A��*�A2�ʱZf��b�2�����JS��7�p���dsXfs����L���b7nc�+��͢�th��:�r�hJa�eH/���"�X[�(W`���>N81�S����
ē	����FF�
��
�.Ɏ����Ɖ6�B�6�����r��DqVJ��&��4O�:�(h� �_f�Y��S��ڑ s|ɝ� 2)
�_��.
��$33+8>�A7�_��k�.B{h��a�pj�╍�L��=f���%��"��)C�f�0+V	�5͖�K��*䣨�,^u��_�N���L�3QfpA�D�s5�%�Y@x��F,�Hvbe��~T�#�P�<��V�M�USU�4$���~��2�1�慱+s�_<$�0�ݟ^�m�#^K[���J���uU�uߋ�C�BDBW��-t<�m
�?�;���(W�q<Vj�G��� ? �'nHЩ�7{��D��z��4�B�2?Y��Y�q:m?R���`雕��a����� r��L��("�g�6=�ﭞ��p��1O������hfT��
��S\
�;���W�N+tR�A�1q!�)�c��N/�H�kvRIT*i��7�>S�����|�������^���ڂ��dW�ؤ(�f�������N,n�� ��ށ{-��{���l5��3�:�y�)�M�{�h�*R^��P�xt`�҄�K$���F��O�� ��G+��y�*�h��C�ΟGc��)���K���7e��f�fi�!���3��$�u�i7�g�|�L8�X�u��v�2�]X��9���pH�$3�m�iAi7��LL����i�E����^�'��:wϭ�A3����M];��Ǳ#�3d |�a(O'۵��֌��Yo��ao���|ݨ<� D�&�����	Ǌ٦pT��T�y7����S��%h�$�1&�s�#���D�^�[��߄M����e.'���E�>7���L�<����U֙�W�mw����Λ�c��ꑢ��x��K�5�����Q9;��B{H	�lџ������X~%��.�"��]=.;nK�FŎf�&W]�
h3�RI��D����{� ���,8�+�Z`q�G��X�<g[���@�-��b�J�b\�7u� gVb4�#:�=R~'�_�k��,��U�c���HO�5���kDY\�?�� �� M4#ug��J9�Q���矌q���_�����VnB��-�1"�?J�c�4�sԁ'埠��{Xr �+l�~����������Yf>\�X���L\��"�h���:Q�<^8�E:;I;���0WeP��E'���/���xC`���e�O�L��ɨ�Zg��(X/����|+,&��~�+��yֳ�7)�.�,��۱��'��8O3|n�?�0I��j�XU�X$~R������9��H^���$
1�9��ɵl�{���u�z��6�	��tel�bRٺ��3kE�O��x6�Ew����
r����E�T��4_�j��>�y�j�'�սoR�J��SF���W���/�8]K)X� 3  U�^���?�w�mv{ʥ��g���=mxW�ۗ�83zz6�{s�A���;A�Ke˰�o����YsK���bE�O��%|�ǔ@r$\{����mSW�
���� eb���v�GK�"WQfLl�˜?{�]���L ŒH�*p�������8�����c�$L�Ҧs-��^��Wk�=���DQ(���uT��
2)���[��7B���	�h��<(��Xb��Y,�.�YxB�	�ˌ�P��fW�_�E������8��\��i�柈�^�����+�`��̭�����n��T������f�e�����;���Y��~���mh�j��2�a@H��6�L�~g���y �eQ�x��oxzQN����v�F[5����'�����C�Ж���NBhm�QPS%|�d-�L��Υ"_W��k�k�y$��\�D���������NS���S�@�Й������K��(���"a����V��kb��e�Sj�Ӑqsцȧ�[������ �Hg�|���#Q���u�C
,"+�ۋ�Y�6�5_�͜]����Bv%e^��\WA���g{v0���U��a�̈́�*.n]� 2r1�Ib1�(X����y��}�82~�'�z��AQT�NY��F��2A�m~쨠ݘ0����Y��O�t� ]Os�/�,x���QJ2{��a�[پ2�S�0���\���J�Ѐ�f'�My��k��_���z�0�1�O;�[Qp_i�<����Ԙ�:u>^˰���ͨ��M����Ƹ}�δ�q�ԑ��RSη[�{����x�E_��'��*x��c��~kۀ��4���ڥfc�����>gj���
J��\6�a�]���;2�SCό0vz?A�Y�����q����G��[��.�C[�C�eX���Wjc5��'@�&��߶È3f����@߉h8[�PϺ?@r���������Tz�O!-��y�ET���ss,Ap�vZ9!t5���>-�'�v��y�o�U;l>*�٧�2�he�'���8�����=�E4�Eu�k'�7����$	�⢽��"�M�K�ޫ��Ie+�Z@���^�ƃx���I�[y-sk����� & Nk��!y`UޠHyl�(�8�Q�&)�2�;U>q��O6�D�澁4�v+�Se��� *��<]��y��w��#��X��p���N#ݎ��d��%�3ݳ�4�{�1���GU��1���B9�r܏yØ!`]���2�0*�p�窙��t]����Dh6➣M���8��D���ugC�¸�%m�.����뗩�aųA;7�]E¨r�VH��%�''��V��{4[���f�T��{�gގ���-��!��Y�R�t>�ͺ�2��0 �;���i	CIEP����Ɩ!ujǌ�.�:���#��$��w����[�^�����5G �l��F�!�~��_f����ݢ�W�D���Z�훱�<���Ѩ?W��;�p.?)��ư�6'q�����>�*0(ȿ>��j+/.a��>yڑ������|���]�IM�iQf�F���
;_1���b%�t޸��9;�4I� !�<.�T��/Qר���~9��]t�r��6֌x����^��R����f,�x�°�i����e�U� �P�.�n� a=%?`>�%f�?C{*��ϙ��Ј���Br1�uKNL�7+^�O��.ϴ����ѭ�(Lm	��ڪ�J���Y$I+X���Š<R�\���m��F��8<��θk�C�k7|�[n��)t�X�9��~�3� ._�0 .,�ڿ�q�W���};�I�gYI�����~{�Z=�;*]eWr��X��˄�1Nn��9�����ۚZg��>ʌya����M��Y9�F���Z�>5�i3�jw�rD�h�}��4���L�!���Z��Rt1x;I�i��U&+�A���~$Q�Xwtg�m�͵J~r�V�ÞD��F�a��u1,�mpj��ax>���{��qh���+�fcW�Rc�����g�x��|��/H%J��$ZJʥݟ�|�2�e�GqFi�B���Z.�-jf0�������DA[��ȏ�J�̰Ӯv+(�bwj<yQǥ��*]�I޺�XO��6_�u��{�\x��!��fg!)$`�)��G��b�j���/^A�P�l��݌���ޯ���`�|�̇[0��ú��AD.�SdI�$6t�cx3�<����ZyљOVEUa�����&�_����N��ufu�fz�w�| �D`8����>��91�G�NoA��9�^`��K�=�IE�]�ރ����=���x�`�ǲG]FMe�o��o���'9��Ο$#1������>������dF�@�6PA�2N�&wՉ.�����{�J|w!�S���zhRՙ^���-8{Ihք��n��������6[��/�ؽNiuI�R�fx�B�K@WRh�(X���\���+#%��
��s�����޽�ޖ�@�ٹ#%t�y UX��c�U��SD�\	��1~�[{�D��n�,3
g�G{0z#g�������N�`BM�"�'K;�L��륌��d�D��*�㳣����{��q_�r��h_)0?��f6��(�av��UD��?v*_�Ͱc8����^$\(ʟ��C���ե߽2/8��<���9�	���	l�
`�K���_x��L��d��J��8��QM�k��,�4��e?Q[���g�;�`D�9�����7�]Y��ߦ����p�U�0P����rҡD���2ܲ�MG�J׭�<' �N�+�\�;�W#�SŤk��J�ǟ8�G��!{ 
�:��ʖ��>(�u3�-Ǜg ��ܯz��֏�.����V~1�4��EAJ��r����*�8Y�L�c�����O����+{J�I���P�F��F��ѪZP��y�����e���G�)�FZU�t�,�����]gS1�%.�ULUr���JU����y�7ѥ�AL�)� a
Bq,�7�������G�$ l���~��*��,Z$H��/��X�#u�1x��d��^��~Z��~\�^]�.��t�"��je� �Q������������	���´v��e��hMP;���Kӗ�]cL�Z���֍f��/WD)!�[�\��\/��h���s	��Ԋ?~!k��O��[h,(�,�Ǜ�~]a��B���Y�	�q�/n
�p,���(�� ��������%tG`�Ե)�E6㡲Zw�������_�^p��#07��FCwd���j-�gO��ٕ͌o��]��XFodom�$��Z1.��m1%��1����2��}���K>��.�q�+�������wU�,�a�av�26Ͳ�n"��Oj��ϋ�oER����3t�Z������@����o�2�� U|��&;���A�~���Ŝ_\<$~1��ᚃ��4�o��΀��c���.����mS=h���"��Z"��W��Օ�T����gG[/bc��I��k�4#䓷/�/+M9"9�����eO�W�p�C���E��ӹ����?Y�)u�)@����aZ�2F�R�С��9��b8Io�n_���	@̇�dM+`���;٠@o:�YL�Χ���Bl�y�s�L�@��B[a^s?y(�jd}R�(�ô�ʇn�N�D/]��K?�Y��� RV��f�9ȧn�HIIQp(��y��������*,��U�B�=2��iY�W��b��ǚ[3�ͽ�K��C��Qkv'\Շ�D3������=�e��� [x�y��6��x�9=���d�1��iu��%�8�&s3�m�FǊ�Aj��]t`~�/5�6N�h��f:�a�>s�*�ʄ��#�-l];R��m�db!�)��
��d ��W{�憖W�~+��xɓ��Ưmb�qؽ�J�o�5� D����a�CKs�$֡�j~�1�ާ��g��L��r/@��)�T��t刚~r�)>mu�k#r:,��f�JJ�����Z��A_��v��B7��[�<\���\�����!l3����}�^���aW����d��T����6���G��H�"���U��]xiᚳ��٠�30�XK��Pl
���(�_�ҹ9��Lͦ(��)Ђ�UyC�s3�8V���y��}��]KL�%C�Bua,S����6 ���|6�D���eS�4����Pqy�$$����d�n�]&y����	�g��F�����?�0D>/r�G�fX��5���m��֐��YC0˦ą2���n��|��)fO@�Q��,�k�"�.
�����?���(K�3XO�ȩ<��OqD*a�sm���:���L���S�r�����0b<.t���T1m�-�y�v�AH�	��.2T��2=	P0������o7��>4���w7{lY��5,3�Ql�����b�=��4Ҹp#�XU�� �T�����U�O��B�ǩ|ew��G�n�Ǚ�4c�A���^聦T^�Y��m�!�&�� ��+�%V���!'�������ǲ6]��;]�=8k�ՖvA?�M�����?!��omp�T�v�Bxq��B��*��ږ�{��`g��H��Q)-O����k�Տ^���!�B$�q�-�q�+u�f~����������J�_û��'qR����};����澋�Ҫ�/W�!h��7Cɡ�Z�X��_��U��ms��.����ᣄ##_�򦁺��~5��� <t�J8B�4��N����qL^�=�2���P#0L�)�s�ֶ��| 1�q�g~�\��;�w��������c4�r��U���
b��J�;�:��U��ǉ�����`$�`��Չ�W��J�Jt]����1q&j���RUw{�8�����e ���.Y=�FJ��m����#����Y�<�6r$�Vy3:���<H�>$*���~��zy7���Z�ד%"_�4o��ɘ�O-��PY-(<���w�T4q#6���_V�*Y���Km|�k�;ϞD��{��A�,Įz1N^z��4.���8D�U[�"j��ȁ!�3�6p�FT�� E{�4t��_��4�?�x���u��j�8��ۡB����xy�ƀ��t�]�3r>��v�>8p.`�8����r4G۵J�%��͍Pk�( (�����*�چ+w I�vl�[s��6�N+LܐO�D �"SAԷF)M��$�(�:t��l��**�^#�CD�?Ї�ԱxùwZlSyzW���ʱ}�C4���� ���Yp��={�H
a��j�N��9�!�/vIΒo�l.����Qy���Ӑ�&z����a����p�X��)N&3C��t�vN�^W�"��&��p���W��ȓ���BY )^���+,��O���`-%K��-E�&���G�א�ܴ���M�MEJ\+�d��0�/�I��em#��	�{���蚆Ϻ�W�1���֊����d\���ۓ�oi�qy�T�U���$��Y�$�C�s+^�XR�6$Q�h4�-�=�=��)�i ���������=Dt}9>�q��L<�r���"�d	;rԸ�%�;�����K����ӵ�c��l���Ŧ���'r�md��+?�:��e��E����n��O}�|L^�_B0�N_$�Մ�|~�jhMK ����i����d�kqk``�5���;T"��)�!��[������s�MD}��3$��Onk#Z��-�@�OK�ݏ� u�)Z;�hRh�-?|+�a����V6�+��'E������V{���Ɉ�#��^����ۦ��2�y$�I�	�Le`����,襄e�	�yy���*LAr�w���&6��ek�\���RUT��-�sf&�^9���������?/9����1˃�i�qE��T�[�Pjh����0�QsxX��J)��i�����@	- �{�(��Wf�I��X�]Q?v�pq%h��%�.M-QP���H���gc~� _z�˛+�mV��@/z����M�3�A�9;g��f�f9�o��3�ɭ�/���DsP �;Z����%� xH��ӂ:z�b0& ��z��C�7B$�y�f�R^��8�}v�/g�*b9z@ A�j.ů�6a����A�rȭ��^n�W�EnV��Sӡ%�O4�U���ΜOICx��
���N���X�G���8ʁ�?����'Bo�s��F3]R�g�_N�'6%�=h�C��o�{�F/AR!��Db��b5�Z��m�G�g{��@�1����.�1D�Y>�����bvq�7�ya-�T)W�����2kGN ����`��>��Ѭ*; ʺN۞f0_�.rn�0����r��x���f�����&j�#Ѩ"ŉc=���L��� ǵt ��(���ý�-WRD6���&�[�%����U=M�Ơ�@��f���B�ʅi+E/|t!��;�6�I���˙B�ش%R<�г8J ��Y�(J���.��7�砟�gz^��5k�3�6���!nw�v����x�X'�0�E��z����a�
�f���M�_��TD��ܘ�����>[����Ys��b3��pE���xJn��� 5��\,t.!}�K[�S���򯻿�݂�74�?%A�R0�����cR0¼���� ')�g)�]ޔ����1�	�3Ij��<�m�PEQ������K��E#EpXI��:8��`�Ӽ�A�����t���V@��͟����c�<s)�z$
iv��;��;��)`��}��(�	ps��Oh�V��	W��;-�Ȑ�n��ߥd�Q׏���F<�gZy�^p���L��WX�J���͈�pb�����/v��kЉ8mq�wp�[������Qs�-������He���qO!@��Ph��
!.����aJ�O���5���A�ޔ�Sڃ�٧�o��Z�C�媢%�W��.�rK
�����m:�h��ᾼ��Sd�MYӲe��Y�g���'�%��b� 4�ʈ��50�-�|�;�/�1� !=Ȃ���q����N{���^��X�
d�Dt'Q)r���>xM㷬�-:�cjxNCȁ�dۈL\���L�`�r�0�]Q%[�a��e$�5��J
�ͺ��S�����&oH8J8�i�z�����S�T3^o347t!5����&A4!`�u��e,-��BI�%+UgϾ�}*��S� Y�����S��e4�2NհlǉRػ]*��l��*q���b���B{O�i�rԸG�2��f�������7�[��46��b�@�xO�tÛ-H�~��U�@��d-K�O(3a���Y��0�\~y�X	v̔bw�[o��17��?�ĳ	�g����b��'i��k��;�?FOZ���-��Q�t4�%	1��O?���ԍ׏D
-|^()�3o �G,ә݅�Ct�@R.�<�=U�RUNH�Fc�1Ie0�jV'钱q?Mբ�J]��4m��z����ʁui]zV�����T'�%��<�y���J�tdi��D�ІP�+rקe\�a�+��4���-T��1gh�P[�o�ltd����v��G�PnZ9�x�f���{�z`@�=��9�]�ΨϪ������'��$�!u��"p�6���"/��1�FD�^�Q$���)7�N`ڛܛ|��>c6�N(��g�o��}�GƻT~����gk�(k�1L۪���}�ƌx_�G���WWd�P��08�X��V�� ��'͹��ȥ�-[F*4�u�c˭���0��
�SUC��+sX�@��Z���p�'�?��Ps����sz�G��_�WIb�ML�= �9�6T��7Λ��΃�)d�|�t25ja��1����r�9h�P�U{�c�̍<�N�(�+���j�֐���/ҕ}��ǉ�eبz���])t���OK|�>y�4:m���!�o�ZJ,���C�7(T�`pS��m���h'�{|�+�l���R	˦Lй��vuׅ�4��73<�e�$�O���ڿٴXA�}��)r�|�y�C���w5"v���þ&<\�N�ۆMՖ4f�߀c3+]F��^���q��̛���%����-a��h���w\}ADϘ#jh�4����z�l��_�tX��RK+��k� a���+KAL�4Z=��C��su��U���6�vd��O��@��vúq�dX23��ǚ��\� �;�`6c4������]]�0b1?W"X��X6]f!�j����w5�cVg�K���s� U�z�����7�5;e�kL��8\�!5�!��s��KԾI�`�9�OQ�0�]+Brxc�.:�qW##���O��Qy7�%�]
zoi���Z��.�O8q�ѐx��ީ���F��{����ԙÄ�)©���n0���7�)�=��1;��]�0�'؉�NI�>�jt	7��M�qQ�&j&cY���Ú�~�������r�*�b0�d�"cBO���D)�f���3�w��u����We�Ò��iy^�x���A��e�O��V��$��s�6�]��ຢ�E�a`I5B �p����?��,����{�.��yo����d�q� �_�����(�G���Ҁ�E�e�5^(\	j��)�x= 0%m-���7q`��Ӂێ�|�)&��pfN�O�� ���D�#ؽJ����D�͘����T�56/�����v�o,�����"RC�\{�0�,�")Qj�#��tWM@��w+��8H-a���mwq@1��)D�����_20���Q��r�U��`Y�$+n9�FәZ��3O�j���6QF��_������F�{~Ҹ���賫"����C�i�ÂG��,��������.���Me��\���u^���q�K\���H�-C'�~n��,�wE
��m'�V�i��[+*�|톭�����X�V��
��������@
-���L�f�ߝ������%�S��Ё�Y�YR�m�9_��=&"�Y͇��wu��qp���`��En�QC���W7d�&Q��?�	g�Y[R�����wU����!"��p_�%R� ���
�ξ����R�T:�Y��b�i�����mГ]Žz��D�	�t�e�#�)S����@3s<G1��ߩ�D�Gu�N)��T&}��kJ#�)և@��8�ҟ�®�4��o����t��q,R=�`q��27�F��������%R����ý��y�l��#&��45K�֐�0��m����d�@��F�Cv,�%�O�<WL]Y���J@]Ok��E�x�����ZI��q�SƠ�>>��S>O��cz��?��{��(9���&��]f�E�fN�b舡3F�� ?O )-LL')oK��~�X�^�4t�A��e�ה���m ��3��XDzLʚĔ�t4������\?
�M���*?��$�?�@����ofI�A�A��}nj�uo�*��f�kS����@���<xF_�CW����|؊9F���Ba���	��A��A�ˣ�,K�2��*{h<�'̮S��љ��"�����C|.�&A~O�V*迣��e�>�O�+K��T��D�l�E�^C�(�zn�\6wɲ�r��Y��Sm�r)� M�Ou�X6T�%�����蜥lm����]n �)��!B�Z`�r�Вһy�gK@�3Q2��� ���P�kF&��FHB��{a�7{=�O7�Z]��,�����d� i} ��/@��6��j�d�J�..��(�B�rC��o{+���&,8Ԣ�@%WM<>��ZP�,kS.]b�3:d�-�Ժ�_˽�v~rb�;���������fe��)/q*(yuYd�Q�rgm��&�i,�����4��b��N/��VN���m�f' �Y����"�Juf��n��.Pl�צּ˪l��4�o�g)u��u#���Rx�;D!�.1R"<����u��B|���u��,景�mMC/��!#>%����:]��V��P_��;5�ɼ�K*z��9�>_L�Q1��$�{v[����^=���]-Jq�����T�-�,��H��H<#����SXY_�����XS��﵇��d���F��_�#�#S�[������YW�ǧ�7�Y�X������y�R�!ͧ����h�#�|��ݜ:8o�c2�U|�.mL�1�C@���X��T�gWz(q7T'"���T�<|D�-��H����O4�R#A�~��2m�!���|���ѹ�L�I�V�吩f�e�r�Q���#�/�+�3㐕�}(���CB�C��I���V���*	u&1��� (R<�أ�m3�e�eyØ��!Z�4��2@=�rvb���w+ɛmW��WgԊ]��2�6%�xTM]�,��=Yq���^C��O���ُ���`��)�ԯ[�Ru�I�SNZ3�
`}褋]�I��~����������艱v����Й3J8��.��f���衫��:<�uI���g��%�N��S<m(��+m5���Uf>qL����R�b����d�6��x�Ԩ�$K{�RF�y���!��%�}� ̊MUp�ܢ:B7����ſJ�P����W5��j�ؚ����>১�Zb�?��zݍ�h9�3bg>祐,0�F��w��D�v��c�ykS�H�7�uSK�W��ʫ�"j��5�p������#*�R�
�Y�gDw���y��z���&��������|x��j�%f������'�,=V4.�e��2�i��b��@�R�J�||�Q��J���LH(�FY����K�{�`aN{쭋|�^:<�QPf��!�1 A�*�/)(t���\gzҺ��u6#�2�Q�
�A�@�'�ߊp�9����t^	k�?��_��\"!�A��� Ȋ�h�CAy_u���8�&����N�N��| ���X|ΒG�]��t�>��t(���t) ���C�c��7ي)_zD�p�^9�)���� B�R,Ov��Ǽ�z��u����Y��ǞuZ��3�hn�{�*֚!�<�G�n4��'Z�A�}!�Aԥ��r�j�x[�@��J8�`K�����i1m=Pa� _b}@��4�Y^8}s�>�cC{m�[z*C�mD�<ԕ������c.�h�-U���\����=>�$� H8?��Ɇ�:�����帴��]������4ë+����3�ư��^�o�!�� y��֍���X�P!ACl���/�v����y8����m�!
F!����lt}�B�R��|&&[��U�n���q���Y��0f�A/3�Od;���z��goдs�z��#�����*��V!3|"��Y���Zu|sL*��o2�@ޟБ�Ju����C�6�|��B��`�I�H{?�R���	�E׭�p����v��"�܂�&�=�eI��:t�ae��Y+l��BEe~�Ԭ�:�	�qN�i���ϛ���$��P�7=*k'�{��_W�k��Zn���frK{ �qy�=�̼TrlQ�P�U�����_��ѡs?�_'|�0�yfIu`4�]��r��|Xw�g�K>̖��*~�2�q"�l~�2���Y?�� ���_X�� ����/�\�'���|���s|b�z�C�ˊ�R(F�Z�1:��'�~�\�f�����t���\�37�M��+/��jK��'��)�0����M��Re�(P���X72�J�	�Z�8��E��w c����2=FA���2M/K*H�y��ƫ��Gh:�bP.U\��C����HBd�i�(�7�l��-�I�s\)�/�c�U!m���s��}=�ǃ��� ���ܢl�.AUiuL2�&Gە�P=?��=��D~B�<�4Z����J�{��_fcnz`�ܗY���"qJ�r��U�G��y�PU�IP���U#�D{����k�Z�]��l@tm%�>&���wEh����M�ɢ�dx^s�7�.H��2Ϛ	�J� �����f7��t�w�wL�d� Ȧ�r��.8MS���#��5���F����Y�
f%]f��9������9��t��s/�����E�
����1nG�|*^{M����v�o���mƼ�R��!w�J��W��zQ>ƩȘ�l�z��.�8�vL�n��,1��bJ�oXԲ��^A�x�Qb(�M���O�i0(g�;Q��=� Ees:no��aRVy�6��9P��lm�v�BLW�P�C]��X�L]�{AvLl�E���Y�7�\���O:7�QQ1�IR��p�����څv�|3e�o)��h_�������#u�ś�~�Z��{���#��Q��G�3jkv;�r+�����Ԑ�r=��"�9g!fgk{���^��Q�\Ė$�"��IBf�h��u|�\�7��OO��������iR�Gb|�4�w��5�cfڱl���z����!M��7{��Z߇T���^0���Ż��|���y�������,�\�
�l�|%����Z��$��#���V�^�T~��uSn�ka�?�L%�ls��d~1�������t�f1Au�]����u�l��U<��k�5���}X�Z� �88%#�C�S�X�cW[����w�5^0Ȇ��)�%�������-���_�T�`s��m��f��d��gq���s���`��A��	_)�l$_iکsi�g�]�٘��~��!�� �b虰�(�ܶΈ�4�L��P��<�lMC�N�o�*��&t����, �>9Y=-o�O�i�RW���"h�ɃW̾��E��G��<Þ�K��B��&�����݅�X�Bx��G43���ID|`9o�
���8����
��0bp!b�ơ���s���uEB�G�� u�p�ֳ�-O,+���6�ߠ�O��|����P���	/��鶆�:�Q ��o��i6��������ܑ�fUw�68�z�"�9D$�S���+G�۪�7Wsj���<�=剄����h�Jab�zlz���d�D��:Hf���'��a��`g![4�R���؉�O�.!�П���XHh�-܎�<���f�!����ې�Gz�	ù'�do5MO2�d)��B�FJ�qsk��>�ѻ���#s��<�Hy�we~�	����c����Jwϟ:.�-�tT�jS��^m�X:*���Cn+����-�*����с~'Z楲+��(ab�[��8&*M>\��R�"��yQ���K�/��yD��5�<���������Y��/?��.�H��?X�p��@�9I�Jp�<��"����}��u��� m|k�U�U%��@?m�V={,�|���K2�0Eg�u��'�V��_B��?�::Z��)]���_��D8��Gj��}�_���˚��5�N�Z��0��t�U�F�Bl4Mޕ��
1�̘���,��,�[Po��Y���|2E�"p`y�G�q	�PD��m���I�p��7r�H����do�*fX|��@�+÷�����f���HXp+~u�I_�	^}|����A&Z"yY63?_�h��v�`vزA�_��M8��wf����ĝz�HzF�~?�B�����}���D@������-]4^Կ�$�n�)��U�k5���T*>ɝ|�5LE<�6�����KG�|X�0'������^��"�InL]�Mjhç楼Gty�l�%t�脑x#(�~�o��(���jF��1<
8zh��e']y�^�h5��7v<�o�܌׿���n�D�V�L��8�x�`�ZDE��j�P�Zע �3��!wx�\Z9u����R��*	%�&�� �0���7��v�Zo�� �r�\��R�]�(���P�}Ҷ2�#@&�R��	�4����A�Eש̬��@��N&/�N��Zm��픱�Dy�W��"O%�OTQx5��k���ju�1�j�&��UM�Ć!�%�����Us�ha�"�S �)����_<Ŏ��1�d�眙���BM�s��<Y�xng��Cu�Г����pe�s���mԊ��ٶi�M�/���t��y)0	���䙍���yl�S�>/�j�^P�O(#�[_Ya��!�<ȽTjL�=�8�m@��P������N���V��g�ߞ�O�
,54o��0��j�$3gN4�p�ݔ<6�	�n�5,�y�P�pbS��	�P�;$*.s���,������Vj�u��Y4��ޠԧ�Ej�{2��)@�g0j��w�>�ٟ�%�\��~�d��x�?�k����i���B�D�ic��;9'�&奈1e]'а �63z��7I	-ԝPV�����a
 ����U��f�i�e$ ��8�I�>�u|��A�)��I��&C�J�Cھ���P�������y
�e�c�/�;�
>�WM�����8�9��؛Y݇eJ�w�\sR����$�Ё5x�'��.@���b&��M�T�� Y�.�ÍS�I�Z����������Ox2	��Ri=;Q�9��eX�z(P6n�n}uqP#�ɧy�x�X3{�#�g	<N6�ɖ���5Է��!F圾���w	u��7�LǕ#N��^����ו�%�_���=(HX�,������rM rF���@�/�K{Έ2r�=� ���;�N:��٘f��p��B٦��2xD��~'6�PYT��lR��v�g�0/��崋sV9J3Q�nsј�k����p��l�wd�I����}k�z&~�7���h��!#�W{]
��RXpI��a����o��}��ٶ�4B=ff�b'�|���da��T�>��k�� 
 8��>�(�dc�0�v6��1��o�K7"��n�e;��g��,��R#
�K1V�ء�I��q#�.W���?n�+ET൙��6�:���D7�-�V4��o�1��%9W�!��Y��Y��P�ʱQa*(���	E��~�6�dr�S���pѢh!o?�2E}t�ʑ<E�8}?��%wh�����]E�N���v�z�$�`*i��,xߗ���s ;a��&��b�Ƶ