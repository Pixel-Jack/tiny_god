// HDMI_QSYS.v

// Generated using ACDS version 13.0 156 at 2018.10.01.16:32:46

`timescale 1 ps / 1 ps
module HDMI_QSYS (
		input  wire       clk_clk,                                  //                               clk.clk
		input  wire       reset_reset_n,                            //                             reset.reset_n
		output wire [7:0] led_external_connection_export,           //           led_external_connection.export
		inout  wire       i2c_sda_external_connection_export,       //       i2c_sda_external_connection.export
		output wire       i2c_scl_external_connection_export,       //       i2c_scl_external_connection.export
		input  wire       hdmi_tx_int_n_external_connection_export  // hdmi_tx_int_n_external_connection.export
	);

	wire         pll_sys_outclk0_clk;                                                                               // pll_sys:outclk_0 -> [addr_router:clk, addr_router_001:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, hdmi_tx_int_n:clk, hdmi_tx_int_n_s1_translator:clk, hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:clk, hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, i2c_scl:clk, i2c_scl_s1_translator:clk, i2c_scl_s1_translator_avalon_universal_slave_0_agent:clk, i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, i2c_sda:clk, i2c_sda_s1_translator:clk, i2c_sda_s1_translator_avalon_universal_slave_0_agent:clk, i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, irq_mapper:clk, jtag_uart:clk, jtag_uart_avalon_jtag_slave_translator:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, led:clk, led_s1_translator:clk, led_s1_translator_avalon_universal_slave_0_agent:clk, led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, limiter:clk, limiter_001:clk, nios2_qsys:clk, nios2_qsys_data_master_translator:clk, nios2_qsys_data_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_instruction_master_translator:clk, nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_jtag_debug_module_translator:clk, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, onchip_memory2:clk, onchip_memory2_s1_translator:clk, onchip_memory2_s1_translator_avalon_universal_slave_0_agent:clk, onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller:clk, sysid_qsys:clock, sysid_qsys_control_slave_translator:clk, sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:clk, sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer:clk, timer_s1_translator:clk, timer_s1_translator_avalon_universal_slave_0_agent:clk, timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk]
	wire         nios2_qsys_instruction_master_waitrequest;                                                         // nios2_qsys_instruction_master_translator:av_waitrequest -> nios2_qsys:i_waitrequest
	wire  [20:0] nios2_qsys_instruction_master_address;                                                             // nios2_qsys:i_address -> nios2_qsys_instruction_master_translator:av_address
	wire         nios2_qsys_instruction_master_read;                                                                // nios2_qsys:i_read -> nios2_qsys_instruction_master_translator:av_read
	wire  [31:0] nios2_qsys_instruction_master_readdata;                                                            // nios2_qsys_instruction_master_translator:av_readdata -> nios2_qsys:i_readdata
	wire         nios2_qsys_instruction_master_readdatavalid;                                                       // nios2_qsys_instruction_master_translator:av_readdatavalid -> nios2_qsys:i_readdatavalid
	wire         nios2_qsys_data_master_waitrequest;                                                                // nios2_qsys_data_master_translator:av_waitrequest -> nios2_qsys:d_waitrequest
	wire  [31:0] nios2_qsys_data_master_writedata;                                                                  // nios2_qsys:d_writedata -> nios2_qsys_data_master_translator:av_writedata
	wire  [20:0] nios2_qsys_data_master_address;                                                                    // nios2_qsys:d_address -> nios2_qsys_data_master_translator:av_address
	wire         nios2_qsys_data_master_write;                                                                      // nios2_qsys:d_write -> nios2_qsys_data_master_translator:av_write
	wire         nios2_qsys_data_master_read;                                                                       // nios2_qsys:d_read -> nios2_qsys_data_master_translator:av_read
	wire  [31:0] nios2_qsys_data_master_readdata;                                                                   // nios2_qsys_data_master_translator:av_readdata -> nios2_qsys:d_readdata
	wire         nios2_qsys_data_master_debugaccess;                                                                // nios2_qsys:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_data_master_translator:av_debugaccess
	wire         nios2_qsys_data_master_readdatavalid;                                                              // nios2_qsys_data_master_translator:av_readdatavalid -> nios2_qsys:d_readdatavalid
	wire   [3:0] nios2_qsys_data_master_byteenable;                                                                 // nios2_qsys:d_byteenable -> nios2_qsys_data_master_translator:av_byteenable
	wire         nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                           // nios2_qsys:jtag_debug_module_waitrequest -> nios2_qsys_jtag_debug_module_translator:av_waitrequest
	wire  [31:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                             // nios2_qsys_jtag_debug_module_translator:av_writedata -> nios2_qsys:jtag_debug_module_writedata
	wire   [8:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address;                               // nios2_qsys_jtag_debug_module_translator:av_address -> nios2_qsys:jtag_debug_module_address
	wire         nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write;                                 // nios2_qsys_jtag_debug_module_translator:av_write -> nios2_qsys:jtag_debug_module_write
	wire         nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_read;                                  // nios2_qsys_jtag_debug_module_translator:av_read -> nios2_qsys:jtag_debug_module_read
	wire  [31:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                              // nios2_qsys:jtag_debug_module_readdata -> nios2_qsys_jtag_debug_module_translator:av_readdata
	wire         nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                           // nios2_qsys_jtag_debug_module_translator:av_debugaccess -> nios2_qsys:jtag_debug_module_debugaccess
	wire   [3:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                            // nios2_qsys_jtag_debug_module_translator:av_byteenable -> nios2_qsys:jtag_debug_module_byteenable
	wire  [31:0] onchip_memory2_s1_translator_avalon_anti_slave_0_writedata;                                        // onchip_memory2_s1_translator:av_writedata -> onchip_memory2:writedata
	wire  [16:0] onchip_memory2_s1_translator_avalon_anti_slave_0_address;                                          // onchip_memory2_s1_translator:av_address -> onchip_memory2:address
	wire         onchip_memory2_s1_translator_avalon_anti_slave_0_chipselect;                                       // onchip_memory2_s1_translator:av_chipselect -> onchip_memory2:chipselect
	wire         onchip_memory2_s1_translator_avalon_anti_slave_0_clken;                                            // onchip_memory2_s1_translator:av_clken -> onchip_memory2:clken
	wire         onchip_memory2_s1_translator_avalon_anti_slave_0_write;                                            // onchip_memory2_s1_translator:av_write -> onchip_memory2:write
	wire  [31:0] onchip_memory2_s1_translator_avalon_anti_slave_0_readdata;                                         // onchip_memory2:readdata -> onchip_memory2_s1_translator:av_readdata
	wire   [3:0] onchip_memory2_s1_translator_avalon_anti_slave_0_byteenable;                                       // onchip_memory2_s1_translator:av_byteenable -> onchip_memory2:byteenable
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                            // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                              // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire   [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                             // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                  // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                   // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                               // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire  [15:0] timer_s1_translator_avalon_anti_slave_0_writedata;                                                 // timer_s1_translator:av_writedata -> timer:writedata
	wire   [2:0] timer_s1_translator_avalon_anti_slave_0_address;                                                   // timer_s1_translator:av_address -> timer:address
	wire         timer_s1_translator_avalon_anti_slave_0_chipselect;                                                // timer_s1_translator:av_chipselect -> timer:chipselect
	wire         timer_s1_translator_avalon_anti_slave_0_write;                                                     // timer_s1_translator:av_write -> timer:write_n
	wire  [15:0] timer_s1_translator_avalon_anti_slave_0_readdata;                                                  // timer:readdata -> timer_s1_translator:av_readdata
	wire   [0:0] sysid_qsys_control_slave_translator_avalon_anti_slave_0_address;                                   // sysid_qsys_control_slave_translator:av_address -> sysid_qsys:address
	wire  [31:0] sysid_qsys_control_slave_translator_avalon_anti_slave_0_readdata;                                  // sysid_qsys:readdata -> sysid_qsys_control_slave_translator:av_readdata
	wire  [31:0] i2c_sda_s1_translator_avalon_anti_slave_0_writedata;                                               // i2c_sda_s1_translator:av_writedata -> i2c_sda:writedata
	wire   [1:0] i2c_sda_s1_translator_avalon_anti_slave_0_address;                                                 // i2c_sda_s1_translator:av_address -> i2c_sda:address
	wire         i2c_sda_s1_translator_avalon_anti_slave_0_chipselect;                                              // i2c_sda_s1_translator:av_chipselect -> i2c_sda:chipselect
	wire         i2c_sda_s1_translator_avalon_anti_slave_0_write;                                                   // i2c_sda_s1_translator:av_write -> i2c_sda:write_n
	wire  [31:0] i2c_sda_s1_translator_avalon_anti_slave_0_readdata;                                                // i2c_sda:readdata -> i2c_sda_s1_translator:av_readdata
	wire  [31:0] i2c_scl_s1_translator_avalon_anti_slave_0_writedata;                                               // i2c_scl_s1_translator:av_writedata -> i2c_scl:writedata
	wire   [1:0] i2c_scl_s1_translator_avalon_anti_slave_0_address;                                                 // i2c_scl_s1_translator:av_address -> i2c_scl:address
	wire         i2c_scl_s1_translator_avalon_anti_slave_0_chipselect;                                              // i2c_scl_s1_translator:av_chipselect -> i2c_scl:chipselect
	wire         i2c_scl_s1_translator_avalon_anti_slave_0_write;                                                   // i2c_scl_s1_translator:av_write -> i2c_scl:write_n
	wire  [31:0] i2c_scl_s1_translator_avalon_anti_slave_0_readdata;                                                // i2c_scl:readdata -> i2c_scl_s1_translator:av_readdata
	wire  [31:0] led_s1_translator_avalon_anti_slave_0_writedata;                                                   // led_s1_translator:av_writedata -> led:writedata
	wire   [1:0] led_s1_translator_avalon_anti_slave_0_address;                                                     // led_s1_translator:av_address -> led:address
	wire         led_s1_translator_avalon_anti_slave_0_chipselect;                                                  // led_s1_translator:av_chipselect -> led:chipselect
	wire         led_s1_translator_avalon_anti_slave_0_write;                                                       // led_s1_translator:av_write -> led:write_n
	wire  [31:0] led_s1_translator_avalon_anti_slave_0_readdata;                                                    // led:readdata -> led_s1_translator:av_readdata
	wire  [31:0] hdmi_tx_int_n_s1_translator_avalon_anti_slave_0_writedata;                                         // hdmi_tx_int_n_s1_translator:av_writedata -> hdmi_tx_int_n:writedata
	wire   [1:0] hdmi_tx_int_n_s1_translator_avalon_anti_slave_0_address;                                           // hdmi_tx_int_n_s1_translator:av_address -> hdmi_tx_int_n:address
	wire         hdmi_tx_int_n_s1_translator_avalon_anti_slave_0_chipselect;                                        // hdmi_tx_int_n_s1_translator:av_chipselect -> hdmi_tx_int_n:chipselect
	wire         hdmi_tx_int_n_s1_translator_avalon_anti_slave_0_write;                                             // hdmi_tx_int_n_s1_translator:av_write -> hdmi_tx_int_n:write_n
	wire  [31:0] hdmi_tx_int_n_s1_translator_avalon_anti_slave_0_readdata;                                          // hdmi_tx_int_n:readdata -> hdmi_tx_int_n_s1_translator:av_readdata
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest;                    // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_instruction_master_translator:uav_waitrequest
	wire   [2:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount;                     // nios2_qsys_instruction_master_translator:uav_burstcount -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata;                      // nios2_qsys_instruction_master_translator:uav_writedata -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [20:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_address;                        // nios2_qsys_instruction_master_translator:uav_address -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock;                           // nios2_qsys_instruction_master_translator:uav_lock -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_write;                          // nios2_qsys_instruction_master_translator:uav_write -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_read;                           // nios2_qsys_instruction_master_translator:uav_read -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata;                       // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_instruction_master_translator:uav_readdata
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess;                    // nios2_qsys_instruction_master_translator:uav_debugaccess -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable;                     // nios2_qsys_instruction_master_translator:uav_byteenable -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid;                  // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_instruction_master_translator:uav_readdatavalid
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest;                           // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_data_master_translator:uav_waitrequest
	wire   [2:0] nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount;                            // nios2_qsys_data_master_translator:uav_burstcount -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_qsys_data_master_translator_avalon_universal_master_0_writedata;                             // nios2_qsys_data_master_translator:uav_writedata -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [20:0] nios2_qsys_data_master_translator_avalon_universal_master_0_address;                               // nios2_qsys_data_master_translator:uav_address -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_lock;                                  // nios2_qsys_data_master_translator:uav_lock -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_write;                                 // nios2_qsys_data_master_translator:uav_write -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_read;                                  // nios2_qsys_data_master_translator:uav_read -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_qsys_data_master_translator_avalon_universal_master_0_readdata;                              // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_data_master_translator:uav_readdata
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess;                           // nios2_qsys_data_master_translator:uav_debugaccess -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable;                            // nios2_qsys_data_master_translator:uav_byteenable -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid;                         // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_data_master_translator:uav_readdatavalid
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // nios2_qsys_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;              // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;               // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_jtag_debug_module_translator:uav_writedata
	wire  [20:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                 // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_jtag_debug_module_translator:uav_address
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                   // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_jtag_debug_module_translator:uav_write
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                    // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_jtag_debug_module_translator:uav_lock
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                    // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_jtag_debug_module_translator:uav_read
	wire  [31:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                // nios2_qsys_jtag_debug_module_translator:uav_readdata -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // nios2_qsys_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;              // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_jtag_debug_module_translator:uav_byteenable
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;            // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [96:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;             // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;            // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [96:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // onchip_memory2_s1_translator:uav_waitrequest -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory2_s1_translator:uav_burstcount
	wire  [31:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory2_s1_translator:uav_writedata
	wire  [20:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory2_s1_translator:uav_address
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory2_s1_translator:uav_write
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory2_s1_translator:uav_lock
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory2_s1_translator:uav_read
	wire  [31:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // onchip_memory2_s1_translator:uav_readdata -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // onchip_memory2_s1_translator:uav_readdatavalid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory2_s1_translator:uav_debugaccess
	wire   [3:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory2_s1_translator:uav_byteenable
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [96:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [96:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire  [20:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                 // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [96:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [96:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // timer_s1_translator:uav_waitrequest -> timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_s1_translator:uav_burstcount
	wire  [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_s1_translator:uav_writedata
	wire  [20:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_s1_translator:uav_address
	wire         timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_s1_translator:uav_write
	wire         timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_s1_translator:uav_lock
	wire         timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_s1_translator:uav_read
	wire  [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // timer_s1_translator:uav_readdata -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // timer_s1_translator:uav_readdatavalid -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_s1_translator:uav_debugaccess
	wire   [3:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_s1_translator:uav_byteenable
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [96:0] timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [96:0] timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // sysid_qsys_control_slave_translator:uav_waitrequest -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_qsys_control_slave_translator:uav_burstcount
	wire  [31:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                   // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_qsys_control_slave_translator:uav_writedata
	wire  [20:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                     // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_qsys_control_slave_translator:uav_address
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                       // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_qsys_control_slave_translator:uav_write
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                        // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_qsys_control_slave_translator:uav_lock
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                        // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_qsys_control_slave_translator:uav_read
	wire  [31:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                    // sysid_qsys_control_slave_translator:uav_readdata -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // sysid_qsys_control_slave_translator:uav_readdatavalid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_qsys_control_slave_translator:uav_debugaccess
	wire   [3:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_qsys_control_slave_translator:uav_byteenable
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [96:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                 // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [96:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // i2c_sda_s1_translator:uav_waitrequest -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> i2c_sda_s1_translator:uav_burstcount
	wire  [31:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> i2c_sda_s1_translator:uav_writedata
	wire  [20:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_address -> i2c_sda_s1_translator:uav_address
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_write -> i2c_sda_s1_translator:uav_write
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_lock -> i2c_sda_s1_translator:uav_lock
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_read -> i2c_sda_s1_translator:uav_read
	wire  [31:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // i2c_sda_s1_translator:uav_readdata -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // i2c_sda_s1_translator:uav_readdatavalid -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> i2c_sda_s1_translator:uav_debugaccess
	wire   [3:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> i2c_sda_s1_translator:uav_byteenable
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [96:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [96:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // i2c_scl_s1_translator:uav_waitrequest -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> i2c_scl_s1_translator:uav_burstcount
	wire  [31:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> i2c_scl_s1_translator:uav_writedata
	wire  [20:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_address -> i2c_scl_s1_translator:uav_address
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_write -> i2c_scl_s1_translator:uav_write
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_lock -> i2c_scl_s1_translator:uav_lock
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_read -> i2c_scl_s1_translator:uav_read
	wire  [31:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // i2c_scl_s1_translator:uav_readdata -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // i2c_scl_s1_translator:uav_readdatavalid -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> i2c_scl_s1_translator:uav_debugaccess
	wire   [3:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> i2c_scl_s1_translator:uav_byteenable
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [96:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [96:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // led_s1_translator:uav_waitrequest -> led_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // led_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_s1_translator:uav_burstcount
	wire  [31:0] led_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // led_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_s1_translator:uav_writedata
	wire  [20:0] led_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // led_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_s1_translator:uav_address
	wire         led_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // led_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_s1_translator:uav_write
	wire         led_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // led_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_s1_translator:uav_lock
	wire         led_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // led_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_s1_translator:uav_read
	wire  [31:0] led_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // led_s1_translator:uav_readdata -> led_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // led_s1_translator:uav_readdatavalid -> led_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // led_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_s1_translator:uav_debugaccess
	wire   [3:0] led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // led_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_s1_translator:uav_byteenable
	wire         led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // led_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // led_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // led_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [96:0] led_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // led_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [96:0] led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // led_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // hdmi_tx_int_n_s1_translator:uav_waitrequest -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hdmi_tx_int_n_s1_translator:uav_burstcount
	wire  [31:0] hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                           // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hdmi_tx_int_n_s1_translator:uav_writedata
	wire  [20:0] hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_address;                             // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:m0_address -> hdmi_tx_int_n_s1_translator:uav_address
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_write;                               // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:m0_write -> hdmi_tx_int_n_s1_translator:uav_write
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hdmi_tx_int_n_s1_translator:uav_lock
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_read;                                // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:m0_read -> hdmi_tx_int_n_s1_translator:uav_read
	wire  [31:0] hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                            // hdmi_tx_int_n_s1_translator:uav_readdata -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // hdmi_tx_int_n_s1_translator:uav_readdatavalid -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hdmi_tx_int_n_s1_translator:uav_debugaccess
	wire   [3:0] hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hdmi_tx_int_n_s1_translator:uav_byteenable
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [96:0] hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                         // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [96:0] hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;           // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                 // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;         // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [95:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                  // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                 // addr_router:sink_ready -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                  // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid;                        // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [95:0] nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data;                         // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready;                        // addr_router_001:sink_ready -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                   // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [95:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                    // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router:sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [95:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_001:sink_ready -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [95:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_002:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [95:0] timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_003:sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                       // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [95:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                        // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router_004:sink_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [95:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_005:sink_ready -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [95:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_006:sink_ready -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // led_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         led_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // led_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // led_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [95:0] led_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // led_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         led_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_007:sink_ready -> led_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rp_valid;                               // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [95:0] hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rp_data;                                // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_008:sink_ready -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                                       // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                             // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                                     // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [95:0] addr_router_src_data;                                                                              // addr_router:src_data -> limiter:cmd_sink_data
	wire   [8:0] addr_router_src_channel;                                                                           // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                             // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                                       // limiter:rsp_src_endofpacket -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                             // limiter:rsp_src_valid -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                                     // limiter:rsp_src_startofpacket -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [95:0] limiter_rsp_src_data;                                                                              // limiter:rsp_src_data -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [8:0] limiter_rsp_src_channel;                                                                           // limiter:rsp_src_channel -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                             // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         addr_router_001_src_endofpacket;                                                                   // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire         addr_router_001_src_valid;                                                                         // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire         addr_router_001_src_startofpacket;                                                                 // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [95:0] addr_router_001_src_data;                                                                          // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire   [8:0] addr_router_001_src_channel;                                                                       // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire         addr_router_001_src_ready;                                                                         // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire         limiter_001_rsp_src_endofpacket;                                                                   // limiter_001:rsp_src_endofpacket -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_001_rsp_src_valid;                                                                         // limiter_001:rsp_src_valid -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_001_rsp_src_startofpacket;                                                                 // limiter_001:rsp_src_startofpacket -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [95:0] limiter_001_rsp_src_data;                                                                          // limiter_001:rsp_src_data -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [8:0] limiter_001_rsp_src_channel;                                                                       // limiter_001:rsp_src_channel -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_001_rsp_src_ready;                                                                         // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire         rst_controller_reset_out_reset;                                                                    // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, hdmi_tx_int_n:reset_n, hdmi_tx_int_n_s1_translator:reset, hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:reset, hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, i2c_scl:reset_n, i2c_scl_s1_translator:reset, i2c_scl_s1_translator_avalon_universal_slave_0_agent:reset, i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, i2c_sda:reset_n, i2c_sda_s1_translator:reset, i2c_sda_s1_translator_avalon_universal_slave_0_agent:reset, i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, irq_mapper:reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led:reset_n, led_s1_translator:reset, led_s1_translator_avalon_universal_slave_0_agent:reset, led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, nios2_qsys:reset_n, nios2_qsys_data_master_translator:reset, nios2_qsys_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_instruction_master_translator:reset, nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_jtag_debug_module_translator:reset, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory2:reset, onchip_memory2_s1_translator:reset, onchip_memory2_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sysid_qsys:reset_n, sysid_qsys_control_slave_translator:reset, sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer:reset_n, timer_s1_translator:reset, timer_s1_translator_avalon_universal_slave_0_agent:reset, timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         rst_controller_001_reset_out_reset;                                                                // rst_controller_001:reset_out -> pll_sys:rst
	wire         cmd_xbar_demux_src0_endofpacket;                                                                   // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                         // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                 // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [95:0] cmd_xbar_demux_src0_data;                                                                          // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [8:0] cmd_xbar_demux_src0_channel;                                                                       // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                         // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                   // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                         // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                 // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [95:0] cmd_xbar_demux_src1_data;                                                                          // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [8:0] cmd_xbar_demux_src1_channel;                                                                       // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                         // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                               // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                     // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                             // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [95:0] cmd_xbar_demux_001_src0_data;                                                                      // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src0_channel;                                                                   // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                     // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                               // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                     // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                             // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [95:0] cmd_xbar_demux_001_src1_data;                                                                      // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src1_channel;                                                                   // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                     // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                               // cmd_xbar_demux_001:src2_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                     // cmd_xbar_demux_001:src2_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                             // cmd_xbar_demux_001:src2_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [95:0] cmd_xbar_demux_001_src2_data;                                                                      // cmd_xbar_demux_001:src2_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_demux_001_src2_channel;                                                                   // cmd_xbar_demux_001:src2_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                               // cmd_xbar_demux_001:src3_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                     // cmd_xbar_demux_001:src3_valid -> timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                             // cmd_xbar_demux_001:src3_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [95:0] cmd_xbar_demux_001_src3_data;                                                                      // cmd_xbar_demux_001:src3_data -> timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_demux_001_src3_channel;                                                                   // cmd_xbar_demux_001:src3_channel -> timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                               // cmd_xbar_demux_001:src4_endofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                     // cmd_xbar_demux_001:src4_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                             // cmd_xbar_demux_001:src4_startofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [95:0] cmd_xbar_demux_001_src4_data;                                                                      // cmd_xbar_demux_001:src4_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_demux_001_src4_channel;                                                                   // cmd_xbar_demux_001:src4_channel -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                               // cmd_xbar_demux_001:src5_endofpacket -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                     // cmd_xbar_demux_001:src5_valid -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                             // cmd_xbar_demux_001:src5_startofpacket -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [95:0] cmd_xbar_demux_001_src5_data;                                                                      // cmd_xbar_demux_001:src5_data -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_demux_001_src5_channel;                                                                   // cmd_xbar_demux_001:src5_channel -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                               // cmd_xbar_demux_001:src6_endofpacket -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                                     // cmd_xbar_demux_001:src6_valid -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                             // cmd_xbar_demux_001:src6_startofpacket -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [95:0] cmd_xbar_demux_001_src6_data;                                                                      // cmd_xbar_demux_001:src6_data -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_demux_001_src6_channel;                                                                   // cmd_xbar_demux_001:src6_channel -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src7_endofpacket;                                                               // cmd_xbar_demux_001:src7_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src7_valid;                                                                     // cmd_xbar_demux_001:src7_valid -> led_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src7_startofpacket;                                                             // cmd_xbar_demux_001:src7_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [95:0] cmd_xbar_demux_001_src7_data;                                                                      // cmd_xbar_demux_001:src7_data -> led_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_demux_001_src7_channel;                                                                   // cmd_xbar_demux_001:src7_channel -> led_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src8_endofpacket;                                                               // cmd_xbar_demux_001:src8_endofpacket -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src8_valid;                                                                     // cmd_xbar_demux_001:src8_valid -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src8_startofpacket;                                                             // cmd_xbar_demux_001:src8_startofpacket -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [95:0] cmd_xbar_demux_001_src8_data;                                                                      // cmd_xbar_demux_001:src8_data -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_demux_001_src8_channel;                                                                   // cmd_xbar_demux_001:src8_channel -> hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                   // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                         // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                 // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [95:0] rsp_xbar_demux_src0_data;                                                                          // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [8:0] rsp_xbar_demux_src0_channel;                                                                       // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                         // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                   // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                         // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                 // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [95:0] rsp_xbar_demux_src1_data;                                                                          // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [8:0] rsp_xbar_demux_src1_channel;                                                                       // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                         // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                               // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                     // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                             // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [95:0] rsp_xbar_demux_001_src0_data;                                                                      // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [8:0] rsp_xbar_demux_001_src0_channel;                                                                   // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                     // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                               // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                     // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                             // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [95:0] rsp_xbar_demux_001_src1_data;                                                                      // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [8:0] rsp_xbar_demux_001_src1_channel;                                                                   // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                     // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                               // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                     // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                             // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [95:0] rsp_xbar_demux_002_src0_data;                                                                      // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_001:sink2_data
	wire   [8:0] rsp_xbar_demux_002_src0_channel;                                                                   // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                     // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                               // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                     // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                             // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [95:0] rsp_xbar_demux_003_src0_data;                                                                      // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire   [8:0] rsp_xbar_demux_003_src0_channel;                                                                   // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                     // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                               // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                     // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                             // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [95:0] rsp_xbar_demux_004_src0_data;                                                                      // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire   [8:0] rsp_xbar_demux_004_src0_channel;                                                                   // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                     // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                               // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                     // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                             // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [95:0] rsp_xbar_demux_005_src0_data;                                                                      // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire   [8:0] rsp_xbar_demux_005_src0_channel;                                                                   // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                     // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                               // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                     // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                             // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [95:0] rsp_xbar_demux_006_src0_data;                                                                      // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire   [8:0] rsp_xbar_demux_006_src0_channel;                                                                   // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                     // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                               // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                                     // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                             // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [95:0] rsp_xbar_demux_007_src0_data;                                                                      // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire   [8:0] rsp_xbar_demux_007_src0_channel;                                                                   // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                                     // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                               // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                                     // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                             // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [95:0] rsp_xbar_demux_008_src0_data;                                                                      // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire   [8:0] rsp_xbar_demux_008_src0_channel;                                                                   // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                                     // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                                       // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                                     // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [95:0] limiter_cmd_src_data;                                                                              // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [8:0] limiter_cmd_src_channel;                                                                           // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                             // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                      // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                            // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                    // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [95:0] rsp_xbar_mux_src_data;                                                                             // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [8:0] rsp_xbar_mux_src_channel;                                                                          // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                            // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         limiter_001_cmd_src_endofpacket;                                                                   // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         limiter_001_cmd_src_startofpacket;                                                                 // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [95:0] limiter_001_cmd_src_data;                                                                          // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire   [8:0] limiter_001_cmd_src_channel;                                                                       // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire         limiter_001_cmd_src_ready;                                                                         // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                  // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                        // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [95:0] rsp_xbar_mux_001_src_data;                                                                         // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire   [8:0] rsp_xbar_mux_001_src_channel;                                                                      // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                        // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                      // cmd_xbar_mux:src_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                            // cmd_xbar_mux:src_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                    // cmd_xbar_mux:src_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [95:0] cmd_xbar_mux_src_data;                                                                             // cmd_xbar_mux:src_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_src_channel;                                                                          // cmd_xbar_mux:src_channel -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                            // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                         // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                               // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                       // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [95:0] id_router_src_data;                                                                                // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [8:0] id_router_src_channel;                                                                             // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                               // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                  // cmd_xbar_mux_001:src_endofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                        // cmd_xbar_mux_001:src_valid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                // cmd_xbar_mux_001:src_startofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [95:0] cmd_xbar_mux_001_src_data;                                                                         // cmd_xbar_mux_001:src_data -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_001_src_channel;                                                                      // cmd_xbar_mux_001:src_channel -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                        // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire         id_router_001_src_endofpacket;                                                                     // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                           // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                   // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [95:0] id_router_001_src_data;                                                                            // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [8:0] id_router_001_src_channel;                                                                         // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                           // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_demux_001_src2_ready;                                                                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src2_ready
	wire         id_router_002_src_endofpacket;                                                                     // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                           // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                   // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [95:0] id_router_002_src_data;                                                                            // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [8:0] id_router_002_src_channel;                                                                         // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                           // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_demux_001_src3_ready;                                                                     // timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire         id_router_003_src_endofpacket;                                                                     // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                           // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                   // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [95:0] id_router_003_src_data;                                                                            // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [8:0] id_router_003_src_channel;                                                                         // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                           // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_demux_001_src4_ready;                                                                     // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire         id_router_004_src_endofpacket;                                                                     // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                           // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                   // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [95:0] id_router_004_src_data;                                                                            // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [8:0] id_router_004_src_channel;                                                                         // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                           // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_demux_001_src5_ready;                                                                     // i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire         id_router_005_src_endofpacket;                                                                     // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                           // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                   // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [95:0] id_router_005_src_data;                                                                            // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [8:0] id_router_005_src_channel;                                                                         // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                           // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_demux_001_src6_ready;                                                                     // i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire         id_router_006_src_endofpacket;                                                                     // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                           // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                   // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [95:0] id_router_006_src_data;                                                                            // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [8:0] id_router_006_src_channel;                                                                         // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                           // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_demux_001_src7_ready;                                                                     // led_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire         id_router_007_src_endofpacket;                                                                     // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         id_router_007_src_valid;                                                                           // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire         id_router_007_src_startofpacket;                                                                   // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [95:0] id_router_007_src_data;                                                                            // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [8:0] id_router_007_src_channel;                                                                         // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire         id_router_007_src_ready;                                                                           // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire         cmd_xbar_demux_001_src8_ready;                                                                     // hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire         id_router_008_src_endofpacket;                                                                     // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         id_router_008_src_valid;                                                                           // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire         id_router_008_src_startofpacket;                                                                   // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [95:0] id_router_008_src_data;                                                                            // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [8:0] id_router_008_src_channel;                                                                         // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire         id_router_008_src_ready;                                                                           // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire   [8:0] limiter_cmd_valid_data;                                                                            // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire   [8:0] limiter_001_cmd_valid_data;                                                                        // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire         irq_mapper_receiver0_irq;                                                                          // timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                          // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                                          // hdmi_tx_int_n:irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios2_qsys_d_irq_irq;                                                                              // irq_mapper:sender_irq -> nios2_qsys:d_irq

	HDMI_QSYS_nios2_qsys nios2_qsys (
		.clk                                   (pll_sys_outclk0_clk),                                                     //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                         //                   reset_n.reset_n
		.d_address                             (nios2_qsys_data_master_address),                                          //               data_master.address
		.d_byteenable                          (nios2_qsys_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (nios2_qsys_data_master_read),                                             //                          .read
		.d_readdata                            (nios2_qsys_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (nios2_qsys_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (nios2_qsys_data_master_write),                                            //                          .write
		.d_writedata                           (nios2_qsys_data_master_writedata),                                        //                          .writedata
		.d_readdatavalid                       (nios2_qsys_data_master_readdatavalid),                                    //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (nios2_qsys_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (nios2_qsys_instruction_master_read),                                      //                          .read
		.i_readdata                            (nios2_qsys_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (nios2_qsys_instruction_master_waitrequest),                               //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_instruction_master_readdatavalid),                             //                          .readdatavalid
		.d_irq                                 (nios2_qsys_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (),                                                                        //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                         // custom_instruction_master.readra
	);

	HDMI_QSYS_onchip_memory2 onchip_memory2 (
		.clk        (pll_sys_outclk0_clk),                                         //   clk1.clk
		.address    (onchip_memory2_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (onchip_memory2_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (onchip_memory2_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (onchip_memory2_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (onchip_memory2_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (onchip_memory2_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory2_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                               // reset1.reset
	);

	HDMI_QSYS_sysid_qsys sysid_qsys (
		.clock    (pll_sys_outclk0_clk),                                              //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                                  //         reset.reset_n
		.readdata (sysid_qsys_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_qsys_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	HDMI_QSYS_timer timer (
		.clk        (pll_sys_outclk0_clk),                                //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    // reset.reset_n
		.address    (timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                            //   irq.irq
	);

	HDMI_QSYS_jtag_uart jtag_uart (
		.clk            (pll_sys_outclk0_clk),                                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                                //               irq.irq
	);

	HDMI_QSYS_i2c_scl i2c_scl (
		.clk        (pll_sys_outclk0_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (i2c_scl_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~i2c_scl_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (i2c_scl_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (i2c_scl_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (i2c_scl_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (i2c_scl_external_connection_export)                    // external_connection.export
	);

	HDMI_QSYS_i2c_sda i2c_sda (
		.clk        (pll_sys_outclk0_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (i2c_sda_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~i2c_sda_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (i2c_sda_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (i2c_sda_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (i2c_sda_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.bidir_port (i2c_sda_external_connection_export)                    // external_connection.export
	);

	HDMI_QSYS_led led (
		.clk        (pll_sys_outclk0_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (led_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)                    // external_connection.export
	);

	HDMI_QSYS_pll_sys pll_sys (
		.refclk   (clk_clk),                            //  refclk.clk
		.rst      (rst_controller_001_reset_out_reset), //   reset.reset
		.outclk_0 (pll_sys_outclk0_clk),                // outclk0.clk
		.locked   ()                                    //  locked.export
	);

	HDMI_QSYS_hdmi_tx_int_n hdmi_tx_int_n (
		.clk        (pll_sys_outclk0_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                            //               reset.reset_n
		.address    (hdmi_tx_int_n_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hdmi_tx_int_n_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hdmi_tx_int_n_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hdmi_tx_int_n_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hdmi_tx_int_n_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (hdmi_tx_int_n_external_connection_export),                   // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                                    //                 irq.irq
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (21),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (21),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_instruction_master_translator (
		.clk                      (pll_sys_outclk0_clk),                                                              //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                   //                     reset.reset
		.uav_address              (nios2_qsys_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_qsys_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_qsys_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_qsys_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_qsys_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (nios2_qsys_instruction_master_read),                                               //                          .read
		.av_readdata              (nios2_qsys_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (nios2_qsys_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                             //               (terminated)
		.av_byteenable            (4'b1111),                                                                          //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                             //               (terminated)
		.av_begintransfer         (1'b0),                                                                             //               (terminated)
		.av_chipselect            (1'b0),                                                                             //               (terminated)
		.av_write                 (1'b0),                                                                             //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                             //               (terminated)
		.av_lock                  (1'b0),                                                                             //               (terminated)
		.av_debugaccess           (1'b0),                                                                             //               (terminated)
		.uav_clken                (),                                                                                 //               (terminated)
		.av_clken                 (1'b1),                                                                             //               (terminated)
		.uav_response             (2'b00),                                                                            //               (terminated)
		.av_response              (),                                                                                 //               (terminated)
		.uav_writeresponserequest (),                                                                                 //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                             //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                             //               (terminated)
		.av_writeresponsevalid    ()                                                                                  //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (21),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (21),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_data_master_translator (
		.clk                      (pll_sys_outclk0_clk),                                                       //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                            //                     reset.reset
		.uav_address              (nios2_qsys_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_qsys_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_qsys_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_qsys_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_qsys_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_qsys_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_qsys_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_qsys_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (nios2_qsys_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (nios2_qsys_data_master_read),                                               //                          .read
		.av_readdata              (nios2_qsys_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (nios2_qsys_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (nios2_qsys_data_master_write),                                              //                          .write
		.av_writedata             (nios2_qsys_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (nios2_qsys_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                      //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                      //               (terminated)
		.av_begintransfer         (1'b0),                                                                      //               (terminated)
		.av_chipselect            (1'b0),                                                                      //               (terminated)
		.av_lock                  (1'b0),                                                                      //               (terminated)
		.uav_clken                (),                                                                          //               (terminated)
		.av_clken                 (1'b1),                                                                      //               (terminated)
		.uav_response             (2'b00),                                                                     //               (terminated)
		.av_response              (),                                                                          //               (terminated)
		.uav_writeresponserequest (),                                                                          //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                      //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                      //               (terminated)
		.av_writeresponsevalid    ()                                                                           //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_qsys_jtag_debug_module_translator (
		.clk                      (pll_sys_outclk0_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                          //                    reset.reset
		.uav_address              (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                                        //              (terminated)
		.av_burstcount            (),                                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                                        //              (terminated)
		.av_lock                  (),                                                                                        //              (terminated)
		.av_chipselect            (),                                                                                        //              (terminated)
		.av_clken                 (),                                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                        //              (terminated)
		.uav_response             (),                                                                                        //              (terminated)
		.av_response              (2'b00),                                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (17),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory2_s1_translator (
		.clk                      (pll_sys_outclk0_clk),                                                          //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                               //                    reset.reset
		.uav_address              (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_memory2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_memory2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_memory2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_memory2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_memory2_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_memory2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_memory2_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                             //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                      (pll_sys_outclk0_clk),                                                                    //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_byteenable            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_s1_translator (
		.clk                      (pll_sys_outclk0_clk),                                                 //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_qsys_control_slave_translator (
		.clk                      (pll_sys_outclk0_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                      //                    reset.reset
		.uav_address              (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sysid_qsys_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (sysid_qsys_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                                    //              (terminated)
		.av_read                  (),                                                                                    //              (terminated)
		.av_writedata             (),                                                                                    //              (terminated)
		.av_begintransfer         (),                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                    //              (terminated)
		.av_burstcount            (),                                                                                    //              (terminated)
		.av_byteenable            (),                                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                    //              (terminated)
		.av_lock                  (),                                                                                    //              (terminated)
		.av_chipselect            (),                                                                                    //              (terminated)
		.av_clken                 (),                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                //              (terminated)
		.av_debugaccess           (),                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                    //              (terminated)
		.uav_response             (),                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) i2c_sda_s1_translator (
		.clk                      (pll_sys_outclk0_clk),                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (i2c_sda_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (i2c_sda_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (i2c_sda_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (i2c_sda_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (i2c_sda_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) i2c_scl_s1_translator (
		.clk                      (pll_sys_outclk0_clk),                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (i2c_scl_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (i2c_scl_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (i2c_scl_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (i2c_scl_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (i2c_scl_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led_s1_translator (
		.clk                      (pll_sys_outclk0_clk),                                               //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                    //                    reset.reset
		.uav_address              (led_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (led_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (led_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (led_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (led_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (led_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (led_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (led_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (led_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                  //              (terminated)
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_burstcount            (),                                                                  //              (terminated)
		.av_byteenable            (),                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                              //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.av_clken                 (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_debugaccess           (),                                                                  //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hdmi_tx_int_n_s1_translator (
		.clk                      (pll_sys_outclk0_clk),                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address              (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (hdmi_tx_int_n_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (hdmi_tx_int_n_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (hdmi_tx_int_n_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (hdmi_tx_int_n_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (hdmi_tx_int_n_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (89),
		.PKT_PROTECTION_L          (87),
		.PKT_BEGIN_BURST           (76),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.PKT_BURST_TYPE_H          (73),
		.PKT_BURST_TYPE_L          (72),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_TRANS_EXCLUSIVE       (62),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (81),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (82),
		.PKT_THREAD_ID_H           (86),
		.PKT_THREAD_ID_L           (86),
		.PKT_CACHE_H               (93),
		.PKT_CACHE_L               (90),
		.PKT_DATA_SIDEBAND_H       (75),
		.PKT_DATA_SIDEBAND_L       (75),
		.PKT_QOS_H                 (77),
		.PKT_QOS_L                 (77),
		.PKT_ADDR_SIDEBAND_H       (74),
		.PKT_ADDR_SIDEBAND_L       (74),
		.PKT_RESPONSE_STATUS_H     (95),
		.PKT_RESPONSE_STATUS_L     (94),
		.ST_DATA_W                 (96),
		.ST_CHANNEL_W              (9),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (pll_sys_outclk0_clk),                                                                       //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.av_address              (nios2_qsys_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_qsys_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_qsys_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_rsp_src_valid),                                                                     //        rp.valid
		.rp_data                 (limiter_rsp_src_data),                                                                      //          .data
		.rp_channel              (limiter_rsp_src_channel),                                                                   //          .channel
		.rp_startofpacket        (limiter_rsp_src_startofpacket),                                                             //          .startofpacket
		.rp_endofpacket          (limiter_rsp_src_endofpacket),                                                               //          .endofpacket
		.rp_ready                (limiter_rsp_src_ready),                                                                     //          .ready
		.av_response             (),                                                                                          // (terminated)
		.av_writeresponserequest (1'b0),                                                                                      // (terminated)
		.av_writeresponsevalid   ()                                                                                           // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (89),
		.PKT_PROTECTION_L          (87),
		.PKT_BEGIN_BURST           (76),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.PKT_BURST_TYPE_H          (73),
		.PKT_BURST_TYPE_L          (72),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_TRANS_EXCLUSIVE       (62),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (81),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (82),
		.PKT_THREAD_ID_H           (86),
		.PKT_THREAD_ID_L           (86),
		.PKT_CACHE_H               (93),
		.PKT_CACHE_L               (90),
		.PKT_DATA_SIDEBAND_H       (75),
		.PKT_DATA_SIDEBAND_L       (75),
		.PKT_QOS_H                 (77),
		.PKT_QOS_L                 (77),
		.PKT_ADDR_SIDEBAND_H       (74),
		.PKT_ADDR_SIDEBAND_L       (74),
		.PKT_RESPONSE_STATUS_H     (95),
		.PKT_RESPONSE_STATUS_L     (94),
		.ST_DATA_W                 (96),
		.ST_CHANNEL_W              (9),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (pll_sys_outclk0_clk),                                                                //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.av_address              (nios2_qsys_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_qsys_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_qsys_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_qsys_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_qsys_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_qsys_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_001_rsp_src_valid),                                                          //        rp.valid
		.rp_data                 (limiter_001_rsp_src_data),                                                           //          .data
		.rp_channel              (limiter_001_rsp_src_channel),                                                        //          .channel
		.rp_startofpacket        (limiter_001_rsp_src_startofpacket),                                                  //          .startofpacket
		.rp_endofpacket          (limiter_001_rsp_src_endofpacket),                                                    //          .endofpacket
		.rp_ready                (limiter_001_rsp_src_ready),                                                          //          .ready
		.av_response             (),                                                                                   // (terminated)
		.av_writeresponserequest (1'b0),                                                                               // (terminated)
		.av_writeresponsevalid   ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (81),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (82),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (89),
		.PKT_PROTECTION_L          (87),
		.PKT_RESPONSE_STATUS_H     (95),
		.PKT_RESPONSE_STATUS_L     (94),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (96),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_sys_outclk0_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                    //       clk_reset.reset
		.m0_address              (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                            //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                            //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                             //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                          //                .channel
		.rf_sink_ready           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (97),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_sys_outclk0_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                    // clk_reset.reset
		.in_data           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                             // (terminated)
		.csr_read          (1'b0),                                                                                              // (terminated)
		.csr_write         (1'b0),                                                                                              // (terminated)
		.csr_readdata      (),                                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                              // (terminated)
		.almost_full_data  (),                                                                                                  // (terminated)
		.almost_empty_data (),                                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                                              // (terminated)
		.out_empty         (),                                                                                                  // (terminated)
		.in_error          (1'b0),                                                                                              // (terminated)
		.out_error         (),                                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                                              // (terminated)
		.out_channel       ()                                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (81),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (82),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (89),
		.PKT_PROTECTION_L          (87),
		.PKT_RESPONSE_STATUS_H     (95),
		.PKT_RESPONSE_STATUS_L     (94),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (96),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_memory2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_sys_outclk0_clk),                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                           //                .channel
		.rf_sink_ready           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (97),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_sys_outclk0_clk),                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (81),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (82),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (89),
		.PKT_PROTECTION_L          (87),
		.PKT_RESPONSE_STATUS_H     (95),
		.PKT_RESPONSE_STATUS_L     (94),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (96),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_sys_outclk0_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src2_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src2_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src2_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src2_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src2_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src2_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (97),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_sys_outclk0_clk),                                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (81),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (82),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (89),
		.PKT_PROTECTION_L          (87),
		.PKT_RESPONSE_STATUS_H     (95),
		.PKT_RESPONSE_STATUS_L     (94),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (96),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_sys_outclk0_clk),                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                               //                .channel
		.rf_sink_ready           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (97),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_sys_outclk0_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (81),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (82),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (89),
		.PKT_PROTECTION_L          (87),
		.PKT_RESPONSE_STATUS_H     (95),
		.PKT_RESPONSE_STATUS_L     (94),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (96),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_sys_outclk0_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                               //                .channel
		.rf_sink_ready           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (97),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_sys_outclk0_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (81),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (82),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (89),
		.PKT_PROTECTION_L          (87),
		.PKT_RESPONSE_STATUS_H     (95),
		.PKT_RESPONSE_STATUS_L     (94),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (96),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) i2c_sda_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_sys_outclk0_clk),                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                 //                .channel
		.rf_sink_ready           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (97),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_sys_outclk0_clk),                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (81),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (82),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (89),
		.PKT_PROTECTION_L          (87),
		.PKT_RESPONSE_STATUS_H     (95),
		.PKT_RESPONSE_STATUS_L     (94),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (96),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) i2c_scl_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_sys_outclk0_clk),                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                 //                .channel
		.rf_sink_ready           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (97),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_sys_outclk0_clk),                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (81),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (82),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (89),
		.PKT_PROTECTION_L          (87),
		.PKT_RESPONSE_STATUS_H     (95),
		.PKT_RESPONSE_STATUS_L     (94),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (96),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) led_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_sys_outclk0_clk),                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (led_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                             //                .channel
		.rf_sink_ready           (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (97),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_sys_outclk0_clk),                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.in_data           (led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (76),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (81),
		.PKT_SRC_ID_L              (78),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (82),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (89),
		.PKT_PROTECTION_L          (87),
		.PKT_RESPONSE_STATUS_H     (95),
		.PKT_RESPONSE_STATUS_L     (94),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (96),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_sys_outclk0_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                       //                .channel
		.rf_sink_ready           (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (97),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_sys_outclk0_clk),                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	HDMI_QSYS_addr_router addr_router (
		.sink_ready         (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_outclk0_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                     //       src.ready
		.src_valid          (addr_router_src_valid),                                                                     //          .valid
		.src_data           (addr_router_src_data),                                                                      //          .data
		.src_channel        (addr_router_src_channel),                                                                   //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                //          .endofpacket
	);

	HDMI_QSYS_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_outclk0_clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                          //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                          //          .valid
		.src_data           (addr_router_001_src_data),                                                           //          .data
		.src_channel        (addr_router_001_src_channel),                                                        //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                     //          .endofpacket
	);

	HDMI_QSYS_id_router id_router (
		.sink_ready         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_outclk0_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                     //       src.ready
		.src_valid          (id_router_src_valid),                                                                     //          .valid
		.src_data           (id_router_src_data),                                                                      //          .data
		.src_channel        (id_router_src_channel),                                                                   //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                //          .endofpacket
	);

	HDMI_QSYS_id_router id_router_001 (
		.sink_ready         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_outclk0_clk),                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                      //       src.ready
		.src_valid          (id_router_001_src_valid),                                                      //          .valid
		.src_data           (id_router_001_src_data),                                                       //          .data
		.src_channel        (id_router_001_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                 //          .endofpacket
	);

	HDMI_QSYS_id_router_002 id_router_002 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_outclk0_clk),                                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                                //       src.ready
		.src_valid          (id_router_002_src_valid),                                                                //          .valid
		.src_data           (id_router_002_src_data),                                                                 //          .data
		.src_channel        (id_router_002_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                           //          .endofpacket
	);

	HDMI_QSYS_id_router_002 id_router_003 (
		.sink_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_outclk0_clk),                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                             //       src.ready
		.src_valid          (id_router_003_src_valid),                                             //          .valid
		.src_data           (id_router_003_src_data),                                              //          .data
		.src_channel        (id_router_003_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                        //          .endofpacket
	);

	HDMI_QSYS_id_router_002 id_router_004 (
		.sink_ready         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_outclk0_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                             //       src.ready
		.src_valid          (id_router_004_src_valid),                                                             //          .valid
		.src_data           (id_router_004_src_data),                                                              //          .data
		.src_channel        (id_router_004_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                        //          .endofpacket
	);

	HDMI_QSYS_id_router_002 id_router_005 (
		.sink_ready         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_outclk0_clk),                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                               //       src.ready
		.src_valid          (id_router_005_src_valid),                                               //          .valid
		.src_data           (id_router_005_src_data),                                                //          .data
		.src_channel        (id_router_005_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                          //          .endofpacket
	);

	HDMI_QSYS_id_router_002 id_router_006 (
		.sink_ready         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_outclk0_clk),                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                               //       src.ready
		.src_valid          (id_router_006_src_valid),                                               //          .valid
		.src_data           (id_router_006_src_data),                                                //          .data
		.src_channel        (id_router_006_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                          //          .endofpacket
	);

	HDMI_QSYS_id_router_002 id_router_007 (
		.sink_ready         (led_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_outclk0_clk),                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                           //       src.ready
		.src_valid          (id_router_007_src_valid),                                           //          .valid
		.src_data           (id_router_007_src_data),                                            //          .data
		.src_channel        (id_router_007_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                      //          .endofpacket
	);

	HDMI_QSYS_id_router_002 id_router_008 (
		.sink_ready         (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hdmi_tx_int_n_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_outclk0_clk),                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                     //       src.ready
		.src_valid          (id_router_008_src_valid),                                                     //          .valid
		.src_data           (id_router_008_src_data),                                                      //          .data
		.src_channel        (id_router_008_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (82),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (96),
		.ST_CHANNEL_W              (9),
		.VALID_WIDTH               (9),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (pll_sys_outclk0_clk),            //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (82),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (96),
		.ST_CHANNEL_W              (9),
		.VALID_WIDTH               (9),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (pll_sys_outclk0_clk),                //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (pll_sys_outclk0_clk),            //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	HDMI_QSYS_cmd_xbar_demux cmd_xbar_demux (
		.clk                (pll_sys_outclk0_clk),               //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)    //           .endofpacket
	);

	HDMI_QSYS_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (pll_sys_outclk0_clk),                   //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_001_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_001_cmd_src_channel),           //           .channel
		.sink_data          (limiter_001_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_001_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_001_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_001_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),   //           .endofpacket
		.src5_ready         (cmd_xbar_demux_001_src5_ready),         //       src5.ready
		.src5_valid         (cmd_xbar_demux_001_src5_valid),         //           .valid
		.src5_data          (cmd_xbar_demux_001_src5_data),          //           .data
		.src5_channel       (cmd_xbar_demux_001_src5_channel),       //           .channel
		.src5_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_001_src5_endofpacket),   //           .endofpacket
		.src6_ready         (cmd_xbar_demux_001_src6_ready),         //       src6.ready
		.src6_valid         (cmd_xbar_demux_001_src6_valid),         //           .valid
		.src6_data          (cmd_xbar_demux_001_src6_data),          //           .data
		.src6_channel       (cmd_xbar_demux_001_src6_channel),       //           .channel
		.src6_startofpacket (cmd_xbar_demux_001_src6_startofpacket), //           .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_001_src6_endofpacket),   //           .endofpacket
		.src7_ready         (cmd_xbar_demux_001_src7_ready),         //       src7.ready
		.src7_valid         (cmd_xbar_demux_001_src7_valid),         //           .valid
		.src7_data          (cmd_xbar_demux_001_src7_data),          //           .data
		.src7_channel       (cmd_xbar_demux_001_src7_channel),       //           .channel
		.src7_startofpacket (cmd_xbar_demux_001_src7_startofpacket), //           .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_001_src7_endofpacket),   //           .endofpacket
		.src8_ready         (cmd_xbar_demux_001_src8_ready),         //       src8.ready
		.src8_valid         (cmd_xbar_demux_001_src8_valid),         //           .valid
		.src8_data          (cmd_xbar_demux_001_src8_data),          //           .data
		.src8_channel       (cmd_xbar_demux_001_src8_channel),       //           .channel
		.src8_startofpacket (cmd_xbar_demux_001_src8_startofpacket), //           .startofpacket
		.src8_endofpacket   (cmd_xbar_demux_001_src8_endofpacket)    //           .endofpacket
	);

	HDMI_QSYS_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (pll_sys_outclk0_clk),                   //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	HDMI_QSYS_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (pll_sys_outclk0_clk),                   //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	HDMI_QSYS_rsp_xbar_demux rsp_xbar_demux (
		.clk                (pll_sys_outclk0_clk),               //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	HDMI_QSYS_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (pll_sys_outclk0_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	HDMI_QSYS_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (pll_sys_outclk0_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	HDMI_QSYS_rsp_xbar_demux_002 rsp_xbar_demux_003 (
		.clk                (pll_sys_outclk0_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	HDMI_QSYS_rsp_xbar_demux_002 rsp_xbar_demux_004 (
		.clk                (pll_sys_outclk0_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	HDMI_QSYS_rsp_xbar_demux_002 rsp_xbar_demux_005 (
		.clk                (pll_sys_outclk0_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	HDMI_QSYS_rsp_xbar_demux_002 rsp_xbar_demux_006 (
		.clk                (pll_sys_outclk0_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	HDMI_QSYS_rsp_xbar_demux_002 rsp_xbar_demux_007 (
		.clk                (pll_sys_outclk0_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	HDMI_QSYS_rsp_xbar_demux_002 rsp_xbar_demux_008 (
		.clk                (pll_sys_outclk0_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	HDMI_QSYS_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (pll_sys_outclk0_clk),                   //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	HDMI_QSYS_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (pll_sys_outclk0_clk),                   //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready         (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready         (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	HDMI_QSYS_irq_mapper irq_mapper (
		.clk           (pll_sys_outclk0_clk),            //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_qsys_d_irq_irq)            //    sender.irq
	);

endmodule
