��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F�)	�ŀ)v�ޑ"^��F��L�> Ó�����M4G�h�.Yv~��f�+�E�9�?���;�Ω0�4��H�;uS%."q��Zd�/�]�+G|��Ԇբ�n�<!�?�a,��5_��=�n�����~t��^}��ٸ�/��eLУvi�i���m�ޮ%G����i�}	�71\&��cq����+�zE��<�`\�L^�e�|�ی�k��=OV�B�v�@�1�^'盾�R��9��'E�򛚤�p�E^΂�Ok��������aG|#�	[m���}�����R��=��ئ4�r-����[�}�x� �|�LW!�c\j��:���ȳ�oi����_v����jqQ�#�d^��Fџ��<0�
)ߪw�B��ֺo\�s)��M�[��	�h_*9o��E_���]��F~�#?ٌp�&�5d1�)G+��� �n���?z!H��x8��U2�#��#T�I�%j=�մ� �Q��9n��C�)��Y���h2�'����lw��9\7�� �9�`�ꌗe��c^E���2;�%�R��� �w�Pk����9���sr~P����u|&��S�-�}	%N��v��	T)%O̘z#i!_ ���*�w�3�Ļ4�L�~�Ǌ���R�o��%!��V��R�����	+ښu�u��a� b� �$ɓ���������G��*�N�
?A}��02��߫w�<s�O������!&v��šc�lA��&���h�"@$��H��r�l�f)��b8�ۘ7c ���|�(<�1��Yh������*�㋽.L��E0pa'E���d�0E�J���G�?�X��$�fxo�#5�P}����,����w��g�VN�V
�#HȎ��U���̏��;Y��c4�p�C��Y9�\v	�5�MX��Ǌ��%�1��9x��X���Zk���j2 �5)e�-oO�P�]�ѐ��n���F�T����
)�@�s��t�P�܆�,\F�Ehi1�������"W�_e�y�ͦ�>>~�/��};�Ӈ�1�GҢ�m�����
 \ n���&��z��e��� ԺU��欀�Iv�˴��D�}!Kdh@����q(6ڮ��X�J&n��$�wݣY�=^'�1/NΖ�o�y�:ϱ���Ï
IL��i$����AI�
�g��i({w)�9��"畠��������dA`��=R�i)��}2"Tm$l)�2ٽ}ɷCf�&�y�K�E���Hi>���z,��ހZ�SqQ��ۘhyZ/��8��'v_JR�~jw1���n����g���{qE��8a��SE�o�u榩������6Y���R���m�{tA�!��N*N�zk��������n�UYy�W����L�����#�w��3�A�R��̮�KsU�H����U_�وo�d�n�1��t&%��U��D G�W/$Rh	�Ƨ��oQhM�6�w��1,�B!|�o���XO[�&�G[:�F�1:���3����ΐʴ��_76Q֋{s����۱�c_�O9j!�4��:����:l��U1y�J�Cм�6����5j�bf�	�fu�i��}yP�2֜:�~��	��Aw@�TeJ�*	��UyG5��Xz����	aby	J�)*��L{?0��s�BO��D�c�2�)�A��W7a�E��} �<�=�p�W�X- t,�k�yT4<dN�R�
x��3Ŭ����h�1!��j��]&��U"��f*�ڎxA���~�J9��~�kfn�W"�!J#D�����u����M�F�.�Q�M� /���)Dn1�;�Hw�'�?Y'��w�������'���\�BW��B��60��;�3<�{9���s��sg�b���pgpPk��a�Y[���#ʔ9��(��W핃��izh+��+���V�W"�`�-{�%��F�sTR�)����f�e�Z�.?���¡GVG��YH�ܣ����p� ��=k�;y���í�x���ȇ�?��Y1na��2s�cZ3^���{1���O��]`?�W	ʽ�x#VʍQ������z�M��&.sib�Z0O	�3��~��߽-���}��=�=�S����`U��O1�$��9��1�������|*v;��aD�ڳ�����Шvdb�ț���i>�xଆ�X|[0�,LI�)ˌZ�����]��e���t�_�kvf;iP��摴��Ǘ�
�@@��F����?e"ݬֻ��n�Q�F�'G��O���� W��a*������f�"��8Ŷ�p�W.�`�0��ya`�r�|ֲ��2<R�:%�i�cb�:5���4F�Sv[�ʫeq�~5�|�I) ���l|9���뛀G����Ϳ�x�\1�
��N�j��^
H|���=�}�H��X�(�=��N<!��,7��Vu��������	F�#k9�p2�4R~��:�%e0�@6�y��.�[����|%q�Hթ:����]�w�, ��l_�N��P.s�n�/�S�B��<���h�=�iu�p�RL��4�n���6��.)���1�-�^]�*v����p�R�;~�Ad��K1=rM�����4c/�tc�Ò2\ęD�C�k�.���֦�9@��o��VǑ�|�_]$(������$FA@XKS�m+���t�Y'�ߥF�甁~�)[�~�Bm,��� �콼/	��{��&��xɶ\
�4
jZ�F��`�E���*}����e$ T6+���#hMu��h|5|�1�L�U�>h,�"�޲�{��g�w.^�X\/�� P
O.�Yg��C� +C}p�
�kp���|K�6��A��q6���^��޾hAn�OC�G���>���2إ�J�J+�ǿ?-��h94��L�%����c�ͺ(R���]�]�Q���0sc�sտe���I�$F�TeL��>�/��ӣ�IpX���g����R�t����eA:m�a�n)�Q}l'(�^s���VҔ-3EC�Bu�"��5���]BW`t�iQb�	��0w���J9ǛK6e-L���n�7�w���C/c8��@��ު%:�t���a�1���WQr��A�kb����\K�0�Y }�q��?��������>W�C[�-���nh� v��$�kt��v��Ym����lRh�?�/%�im�_�8?E!��%w�]A۱�9�~|;�� �����iZ�,C�X������М�W'�.;�7�������z[�|��r�B}�ǈA�V/ǰ�M:	2���� ��I��piKlI��S4f�� �"���=�>����hj�t��K���xx��L��ko@^�U�ܛ���~���9GF�t�j*ŵ84���Uodp"D��X�Cxɞ>Ql��8�zI��ƿ���x'��^H2���2�X���)�����i��#�7��>H��~���)
P0��h�؄�z"Y�s�ݕGxw���g�yc�X��ͣ$�,'ڍp�V��zRg_J(�!�3{~5��O��D�
�٠��-���P�Dl�����}t�y8Mw޼)��N(l�\�����,~�<EHW��-�(!�a_)FA���i�
2�����P:/i�n��Dd�%�7��\6������W�#F՘քD�y���}�Ka�O�����Mz���O����h �Vn�W���9
������ x(����<����|?������`Z�&8�X�<�V�l����Ν֗�؜��r�g��@e⩉zUI����Tw*>;���3b��;+|;b�UNE� ��APN��)���Xa�9�5Dֽ
vEV������ ������Qm�qι���qU�h���@�����<��cQK���Vj+-[��� � <6Q�K�ω'=P�p�G
PB�E�r�x��o���4��K�ű���? W"�/H4|�w6�KC�ǰj7��ڜȵ(���w��%�����c��8
���w��F��������p�T�(���*=s��ٌ����ӇH8{�"o%'�Uf��@�̣����.CE`�V�@���K��Jo�@0+��%2�}#dف�{��]	8JDnj,����l��{�2,86�z58x
&N4������|��$þA���+�����Xe���6$�P��8T��6�X�{R��h3űi�bj_�T6�gÑ�H���p�r���^�㫼��L��@W2�W�T��
"8�H����~h��x#�aNf���!�����]���@zg��@�puF�5XN-	��!R߁wKb8�T+���MX�$� ��SJkG��w!H�=[?�� �cqc��^��:����?.50ߥF&���Q�I�u�X�Yj�g���G)���Y��hҝ%q����ܯ�t����%�O:|��И}"��Pb=N�,�n@1Ex��8C1�F6��|�(;\��kL�9C��B�)�+���mkҞX/�t��5�ҝTf�jA�2����D����i�o�:B��ƶ���~t:�O�@�9j_A�_���591 �51o��nip{3����M����]ɹR�	���6WR/5��F5�W�8*����"�,��6V��Z	�R�2>�"�\U�K�(��E��o��4jP��X"�i�):d�hqU�>���O��r�F�\��Sf��Y�`�S
Z��C�n��DB.�����?���|V�_�� p���!�7��B���O�x��}W����-��:�p�K6�������0�	�6�.���\���$��Bb���sߩ�-	W��*��:l�zн��Zy�x/�A�W���O�RgW�91��%7M�̮�M�BE�'�8��Y0&�@5﨓��b�T��+!Rw�}�æ9��Z2v��ٺ)�p����R;_I���鼉�������0j������3�2%/�Q$���	Q�)�IƬQ��InZ� �Ј�A&G��q�ɹo��&v�0v�Dmw��X�E��&�i�vT_?�VNW%E�]��Tʊ��I���!���;�:����c�G�D��Јx�n��re&����cLm*���P9��1��RV)��hڶ�����"��xHW)ެ��G]b�S�$Y0��5)���=�av�~��S�:r}+_�C&��*_��!w-O�"u��&g�JW'L�2`5���	��ӽZQv�©%������ 4.�Xznd?H��踉n�o�}udz��E#_�	]"��ju���R�卹�ހ$�V�iv�gyN�珱@��g���h�`�#I�������-���������co���&O�I���3�Y
�!�y)r�X����c�W�ᢁ���x{p��[?o�˗�9OA:�X�8%O)XZ���K�p�L�bH��j�۷!ŕ�&�B|�F�f#�mśE�r��`��dR�s��9�kK�F;2;�7�8׬�v~�#F �=�1�$��UӇ�(�I������a]Q���T������!w:�9g�n�z�-�w}}�<�$��_^��_ЮM4qA��f�Ϧ�$q�u�Ġ��Оˬ6�����c*5�4	�R7'�����F��wf��c�Q��p�F�pF��i�>�b�}��,w�B����4�"h��CbH��t��>�� 1o&��4�1H��F��K%�m�&��fۏ����(�e�1T�s�P�(|*�W/�m�$�nϢ��G��K�?Z���2�00�8n�6�)�x0DW�To :��z>qH���g~tsQ���Wv�+W?RN�0A)^lҟ^������_��{����7*���w�5HO�ħ�.��ߟm r2�
<�8"�E�c���ێ钸 ����X��e$~��;��gͺ�f�_9mStC�n���$��Gd]o��Yq�)0����_��h���qfcE��Ү͑6lZ�|V�j�l�=aR����B�J~YĤ��@�,j.x(�c	����z}s�G��Fy���лf����T�ݦ�@P�@���R��f��/��J��׽��<aCX>~�5��KUDn�t��$���F�%���V2!C��oKȄ\	S�f��	��* -%�=9�x��b���/�Y "];IM�U_���˭y,����v�lR���T�3���M|���2]���
�����˘,{��r߰3n��6�h
���@C�=�J��U��Z�t]mI��3"G��C���);�x�PI�PS�Va���c��g����E���5`.Qky�y�Di���̍qF��x��2ng�$��[�t����%�z�&���cR��nnD�-����V�x)EX)p۔s'@�d��csRq)��jj��ʁlkN�ׅ�����x�(rg`)����h�o��@�v����u��a(d�fL	��Wt�I��"���B��;��NP��W0��qk(Il0��}E�K�إ�ߓ*�����e��Na`=2.OC^�j��.'�񋼂�����;��TU�U/�Y�0|Q,�=
F&ue������L�e�y�@���h4��#Uh$N��Z�������T�6$��_-�Q���X�:���<�wZ|$N�B�x�W��y1��ڣ'�R�uk�Hu3���3A?]�z��S��T��$Z�*�;L?0i�$�\�֕��e�X��� }�k/E�_�[Q[�����5�k-w��rEB��.n
9�>=	3g�N�`>-���FJ��P��%�=�6�.[�g΂��¬}��eJ�4�����V�^!�x�f��p����,�Y�a���Q�cık��6�?��H/Aa
����L���!��F"�Y4����?��N'��q#�H��ev�����4C�9�\��/��Ԇ/�9��eq�F��j13_QpL׸�M�@���4�{�d�)ivr���e2�;�E�g=�	�K��h�ˬB����p���[��m���wF�8,dw�M�;h�� ]��L�Ӽ]��Y�V�am:�������g��9q�����"@�0�[�rY>���e��m6�5	ӵ (n�T��:W'�S�%w<�ڼҴ�r��V[�<ZkV�ky���G�0���H����8p˴P��=�J����!��K���Q�6��q ���cdG�1ǹ�d��aFs�5���J�x�FM�jSߦ�X�<s�j8��z9\��p��-�^
��-K�X�T-�>�.>�g2�i�B�#ou��a� '�;�l�L��\��A���Gp=�uٛw���,����W�*��F��tѤ\K�HoN�XH+�cr����h����/z��$���QU�n�P�H���:�H�e]y�>�:���SXbE1	��k���X�4��Z$� � L���M���d=�������_/JF(M��F/&v5�`�������O�����[�ú ��jk�����t@S�ä�w���ݥ(��6�p�8W��.�Wx��м�u��G�c��/�'z ʍ0`�`i�4E���B�]��r��tnm�"}H߀]��{{ �d��k'���l�+�+��VH$8z��~jY�t��Z�뵎��wF�x��dz�3�k�K��c|���t��iT�� ��?���1Vv"L�����G� 5[w������x��½PX��������n������%r�V�d�
��@A@��u^U|�wV��-�3-<J�j��HK�e��̸tk�Yy���w��!˴�Q�ʽ�6[�o֪�3�?Gud��V~�c	�9Zo6�8�7[x19����nYH��}u2|p��^Bd�˟���	��������g�ݡ6��J�b[0c�X�<�mWS?�g��Yp�N��VH:"���
Ef�Fp�<Hn��CZ��>�y_���8�I���23Zy��B��kF���b$�7�xҬ��B�v�K�h~�Sp࠷�Sf�C5 ��$9��r�o��P��ڭ�'���U6�16�W!+����#Ē6�ڏ�%���rי�E9��ïDgO�sl`�G��YZ���xV}���d���X�p�S�3��Ł�&�b��Ð�:k�Y5���w^eh���پ��H=��o'�}��&)FX����	
��;�)�M=V�M�����{��F[?�iQ�����!�w�	B��� )՜,�=�MH1'ɐ�6�6���[:�G�).��C�_x�oF�7--�!�Ӝ	U>c�3�Z^��`�@��=�s�2Km!l�<�pPP����_��2�#�=gU�a<?��Կ5A'մ�]}߲�Z���a6�L	���'�<��vӅ�2��f  �܊.h�cL�=��ð>����i�ڟY��]6	�ؾ\4�ʻ��9/@�e~ ���C�>7��eF� �-0 ҬաB}=R�>���̵��4 ��I�I��|�)��	����+`���$XB�#�y{1=��&����{el��e֢v�>:{��՛����G����6�|���O|ڰ��gI����}M�jJ��e,uĶ��:�����;ׇ?�w����v�d{g����͙�����IN�� sc��e�|������_��#�r�Ǫ��`���p80$��X�۩F�QtPM�xγ��<�{䙬0����O�(��0�c�l��-�����f-GM�!�4T���n��
4��2�\`W�Ლ��z���'��S��t�9h{u��j�U'������k\?�##1-8�3�ن�4-��ul�3h@��͊
���ȶS�4��1�?pDJ�h嘊��׮�?琯r$hABB؇�W�`��h`2`@��ʴh�Μ�>iGxm�HT<$b�#�N��F�8~,�G�h����8KW'�ƃ�ȸ/P����X�b�A�=�Tk�Pm=��N���bn�tf��	�HGȻ���ܻ��4$zdU���u�v�-���;��U�I��Ю|�Z�3�u+����Cs�n��V5��=��� ������WIC������omF�"�ɬf�x�1+kZ>:�]@��K)�j^�Flj��G�-Fg�S���t����� ���@�(�A ��X��!e���ڹ���x�7�l���w�qhG��U��+�Y'���W��1-�C��]t��������D*8P���]l�E-b�R�海���;d{I��A��AnݿhK6*�&������gg���uů����֓V{��Y�[���sv��R~EO�=�Ŕ��T#[�F��T�N?��F�k�kJf�=�У?jY����R��U�ܾI{�:Q�u�cZ���A}:kD\c?��?!���y�m�{�@\�;n����1={���9��6!<�E�BSU�t+9���@P�:�ӆ��1*��1_=	;���Y��lZ�!j�i'���pX&�W��vsD�m�US� �V�Q|)��Bsm�.��@���g�%���f�9�7O���+py�t>�_������|y�ܒf-k"�PY(S�&�-���D�r0�T�/��1�'X������P��˧
��������mP�%Fa0����9�U����c�w�ܸ2��p��2��T[�W�I�A(/;�_Q���6̥94���V�$}3��@�S��CiۘN��� �!1�ԠRl��:�<΂����c!��9��#U��_,�#QI_ߵ��yÈ�w�xPG���,��lR���f�1���=3�7��| �q�����5�N-J��!ӽZ��L��]8�����a�}޼���6�ǘ�6�x��
#U�?��h���dAaJ��w�W`[��j�ff~�x�_A:��M�0�"�e>}{�W|*�����G��iL� �% ���T��V֠��D09�F�1'ˑ�,c��<����m��٢+[?I��8��ŬV���=�A]K�x�{<��(�g�t��.��ʬ��7��=�M.�I�(�+v��೨���l��A� �(�� .���6�;H1?&�yJ�V�����eVw�Ӓ���կ9����l�!鑵���z\���6,W�q��/�y�m��d��!�|U�	����R�z��	8J.:Q�����S�VZ^X���⦒���[s����ߙa���SJ �Q��]*L��SC�4���}���Ф��V�r�+,�*˫7:���"|� �K�Ə��G>ӳ�Gլ��]t�5�T�'��a�Q��M�WǍ<�9=_I��x��1f�^�
k������n��)�?'���ir�(Cħ�r;����;�Z+%�ͤ�,������A�@��E4"�_�A��?u�g��K�B�O��@����ib��{�F�1o��xd ��2�
�~� �~�{�0����d����������k��7�Ȗp���i�(��Vҽ5�ұ�aP-��q�vt��f�߶���(���M����A��N� ��C���)�=-+|'�Wg�m����rM�S�-i�֩�'��7���oB鄀>����*�{��]ᒻ�'N�;�C�6fg�����B�B�s�B������d�!�����L��4�8O���p����O�����@p�F4��1Z��.�ޏM�-+��!=/,)�����Z7����&ڗC��B�<�t��u�YY�������ț�16SB��߼�����(Oz,vΠ�U]g�H���d�2���?:�1s�����K'���SI:ANj|��+sA���m��Xػm� �0�!��0�C/�2q�)֜̎aK�9������?K|�����O|#�@C���u=B=�{sY�~*^��n�ԁ�z��ى�z�0G���ZNo�h+��Ѡs�u���K��_=T���7�9";���a�$:ڙ�t0h}*9CW��=��x��$���^��Sm`���}���Oè�*>����ע$�rA��yn�W�ƍ�r�*�(�YFr!�-Q_��E�AUuԱ��f�';p�C�BR_�lx�-��"D1� �����w*݋�_�Uc�g���!��_>6&�X���М+���LR�d�zQ ��F���v9HK��1�o���DT,�e� x�VOٿ!a3ʱ{@���
�hT�!_�Ʌ�Ǿ��5� eNy�6/
�j Q��J��P1m,��C���F�:��B��(����Zv��"�]J	x
�p�e�Ԋ�
�����d�"�`��}�>��6ꀃ�3?�I�f~���)��B�W
�{�i����W2�_�)��*~jP8d~Nj��g��jT��j��!�	I3���7�/%{�Il��yWW��s\ ���խw�Wa�����v��y4���~�B����7ב&ɡO[��O-n����.���i��e�Z���Q��a~,G�#�n���.)�Յ?%~W�RH}�����ƪ��2�x�=W��-� I8�^5�#��t�Έ���{���j���F2�x��vϮ�J���͠C�n�T;��D��A٩��ǣ�|�Y���ϼ懊�w�9�����G+��a#�P�8X-�-J�*̗~1_U�aĈ'��H��9�#!<|�{DO�o�o�om�R��������=Rl�O���CӨ�ܤ[ca ���Ǆ :"���/�9S�B�D������yc��V�G�u�b������lq��=��EP�Z8�������X�V[��s���P%��f�w	�[S�m�(I��i�j�U(>4w�ЀV���I��؈m�XK`���X�ȕ)��'g�G�p�U7����IT�������>���JYJ���XߩC�~�fԉ��+�	#����ֱG�pb�Xi���L�Z 7�PK�%&���x��o�(ٍ�����^�9��cd�dO�z�?W���6����bI���#V\�A���2�&t���Mޓٮ��{: ,T�{�ۮ產!0�c�	&Ii��K���;"[��_����˂W�Mu�͈�Bd��а��hU�ͧ[�7�� �{�g݂����\e|�S�~ל�HY�*���e���XM_.�~Q�	��d`X�
*�*�L(�5�)��n�����T������"7#�؈On6Kޑ/�=��3~5��ܔ��'٨��j�rW�3&��@�G*�.��5�[�@��֏}��\T����#ۣ��]�&�⏿܌��5�0�]me��B8��9��=��6r���o�6~�^�z�J��y��`{HO��J�8����됃��&8\\��.�Z�F�;�ܥG0=0_��~�*�^�xc)�1>�iGT��R��غ�^��n�k��������2��L�2�7�N8��i���2mg���q��,v��S���V]Tqd���f嗣X�p�({��4JУ|,�h$+�J�ꩯ��b@�Ok��<�L�����:Ԙ��71Su2���J����U��z��5Ƅ�1An����KI��(y��2�P�� �ƒ�z�QVϩ�����@���z��"�E3�f���a=��CÛA?V�	��*���-��P��뿠�Oih�ai���s�ҩ�ds��V��R}�@J?u�5�����;>�aib=���{���c�&5�1�>_�݅+�ԡ��?��p�(�x�LY|�u��ڧ�a�à�|�[0J�+ZBtQ7�v��?�t|��IV��o��Kb��b�u<g]�5"	^���wy���G�K�w}$t���Ӊ\�Ec1*�}c�6�! ֲ�9N2U� &�.g��f���������� ��O������ﵬ�7��7�<�9�����Qs�O�����dz�]�h�a-�<{�㿷����v$T�F�h< L(���,RVz0.��pe���[V�Y�I�&�N�I��)eIa��A�@}�j�A�����v �h�2�W��_�F�C��j�$!����}�D?�\4���4��U`E]7����E�\��W�F�6�&1��Y�+K�n��B0���0�	�2�S�S��a��	E���G?͕�C	Ⲹ�aa����N�q��]tT�>'�@�l��]�R���w�f���BG(7�"�*�*b�1������%(�4O7o�t�2������F�LA,�^�t����g#A¢:v{�χ?r�M�$��!���n���If���a�gC��;��!��Ar_�i3M�������&��m�եF�'b3����//�U=�����������$�{�A�K:���LE	Hw�ڕ
+-C>x~��F���\Y�y��4ۛ�!�ڊ?��'�+b�� ?(o���tY"ϙ�A�m���L&%��߸\�t��z^�.j��B�üO���_ ��M�~��Sr~�e29r�!7(G��Pv;aYd&m�E�������z�5=�H{^n�k&�F���ߡ�.�"t-H�� `H�)�ַ�&�-�}��N�ޢ[�?��>��z1J��۰^	��U�k�x�ǡf���0�s���[f�rh�8q7�����j�Sc�!L��GO�I+�>��B��6a!�/�L{s;%(/������<G
����c�@V̎�i�,�Z�r˪��?�u*��LC�j8��5��E���ϕ>k
)�Dg.6!ש 8�C���F�a�#�!NJ^�橐'�z)^���eNFOK!.���Z��9iղP����ֿĤ�6�V�rEd�Q����tv��/C�e-��𹹎m�hr��"~�V�������B���K7�����< =;[���>�.�=��\P����P�fҜ��^��o ��N,D5{�>�HZ꫏RvJ/��8�,*�����JB�ȼ?�;���)g��m!�P�:�	"��eM�1�"�Hgq�q�?]�	H&��FC��o���č��p7Mo�jvwB5M�֍1�b������-!��0�b��\x>������[��*�z��oT��+�׵�, Ü؝]���v��La�2���3mͩ3��o�������GCbl� 2����:ƦY���0�������g������}���n��	��h�&��-�#�A�e��q?���{�~wۋ��{}7����,��� a�$���kI��B�$��E��&CN/x<��Z�+��Ծl5y�{���\*^�c�rQ�rw�+��q|�+��!����z��w��C����I�#�t�]*�6���9]w�������C��6�?B��:I��k:Y^����dCW�,i3+^�
ۻ@%������?H�}���ںk�pxB�?<��� s�F��D-m��L_��?`���D2��4'J`;��o�w}��|q��j��.�C�8�E��/ka��vB|�9j�����mX�f���Ae��z�wۼ����15R�H;�]ܾPG�AN��i��PNkx��8i��Ǆ �J�w�@ڦ��%K�67Z�����l�Z�q,��n�1�Q�̐)�W��K�52��d���_|���9����+��%������*�?��s�H���it|Qv�J�i�9���]e�����o��.o�K0<3���S�����d���2i{��dow�ӓe*+vy�A�d�x�i{�l1ͅ�s
3�X��*�l3N8���X��(e���9����E�b8˽��{�O�&tѤ�s엪4
Q�CU�Y!���Qp�`B�V�=�س,�G|�� �#݌�&�T�������t��@݌X��膔��Ԑ�Ͳ-W�̇	��C���2F�>��ZN츥�C�?��ڊ�s���A�C�tr4�̝qc�  0P�e�CFz��G"�
Z�i��0x�$�gW��Of�q+ʂ��� �I)`1�YܕB̲Z�h��^̽w�ə��Լ�},І�,;��1oc��ߑ�1\$k����[<�	��gm�=5Y;� ^�"e&��W��/��@:d,���zJu�w�0諃������3���uu�H�(ı�.=�_��TX�Q廱���aXNU/c�Ie;52X��A��"{n���ZQ�ƻ��������s�,��$^�@$jJ��ka/�6�xl�0<l���Qk������k�m��us��fu�Li��#x���뛂-�g~�f^N
��efl�"3��@p�Q�Z|F��0Q�C�����zap�@�E�Sk��mcfZ��o��.'��{�0��f�`�I��EV�v��]�oS����� 7�3ޮIWkn	�J�Pւ�)�I_)��qv���.���`S�@��4��Z�&���� lh"�u]Ļn8��a
��L�x.��˩ oK���a6�|-d�f�֋v�_~�S�̚�)ڵ]I� ��_����N;#0�����V�^��@�g1��R~�y�5.m�<��DM���=I �S*����f%DE8dk���-"�� 
��9̺%,� �7�� p���u�ã9������"�[�Z) N�����
<�W#-U��μE�i�,���z�搿�嗊�GLr����r�|��je���[>�^�I����0.�v�GQM�od��13�-`��h���lw��{u��������"��c��G��yY�L,���H�� x	E׿�}��a�M�]S����T�c��YȐvj�XЩh4��c�tuʡ���}����y0�����h�����X���s�tg��I���QE1�B��,����
ӱ^��x�n�,�Vh�@%d�
�Ggc�a {�UdM2O�h+J�o����K������E�O��.h�NE�b�T��ɹ�.�
i�'K�K���GJ�%����<��Gl/#�����Z�Q`�����?g�������&\�xN����?,+�&h{�ْǀ��ۏGYE���}��ꂼ;�/�0�ƆE8��o��-�X�N�>����]�R۬<bv9|j�*���oR�2D��lqtZk
�������Ah�(��JK`�����J�[O����
���*�����/��د
��'�⺑Z��ȝ�{(��㱔������V2m���laǚ���W���?Tp�)N}iXA�!M�͚T�ׯ+|
�S�u�&�s����2K��2k/{+?0�dkx���-�n�(��n^.������~�[Ѩ�;-���T?�'�K��+�t�y�.s)��]*&� Fs0{P8��i[N��_���g�h�@@J+�4 e������aZ����u��R����v�2uB^:�|DC�|�����iJ}��O�q4�,�&�]��������9Fa�`@��;�]�m��'8Gؾw*OM�x0>�W���V�J�����*ק�U3���Pl:��!�x�y���(��A�J)��(�2G�ԥ
T�̬���?F�&�Ww��3��7[�II^��Pz�!��ɇ��8��6D��.ʴLQ���+.+��x�c�)d��_Q� �ȍ<��-1 �~��2�`�}["'�9��<�	�[\�E��T�.��3�9k�i{���!��cY_���W����֊~�ANg��f�Tೣ�T�6J��̫MUn����|�1sml�{͒�4>?@���6���&���d%j��R% �R���Ż�J,x�L�>�J;%�4
���JZv�Q}$ �y��N�G�sޣ0��uU���S����F/���T3��dQ��,@�JȆ����"����B��y��l���2�8ȄV��F.@)ߍ���}��X]{&��y r�73˘�f�1W&Oo-�/���X�x
3q̢EI~�t�+ݣҒ�T�&�g�"T����d�����f�t�8>ϑ^%1Q�H"��:?�o�~o_��\����������"Q�.](Y/n�o�U�+������/��Rp��.�)�:��MC�����p�P��@�6�#��98x(so���5�5@�	���9���}��q�Y��{6���^�4��R��ΞL�u�a!�
�]5rT� ��R�{h�BF$�μ&^���K��, ���C�"���7{
T����3�yh������$�L:ߒ�3��v-���x�:�U+6�Yɴ�v(i��R�ofQGO7C���Qs���K̟	7ݶk�-�%%��r�w�18�v}��4�6�f�i��'�z0��b�XM�����,U	��zu%oDA���+�[�TE�%)g�'cZdE�R)�r^9�b�����g�H�0̛�������|�`��V6��4kN	&]���h�����;�|�(�Ӑ,�x��< �^QYe<��n&�#W��L����h�/�ŵ����u`֬�u^1�8u���w�aE''�ax�4�>.�f�{�n���0�.��h�~9�)q�%�no���dG�������=Ơ��.�N������G�����>)@y����革q���pU�[n:[��r�#c�@�i8�	���5m�ƃ�{��;��>c�lOq�P��O)�$R��1����|5�/��
OA��sDBj��x�uώ`�m���@����i����v��l7V���XHLS�~�][D�C��ddHE��������GG1Y��\2.o��1h�Ii�p��/�)�G����|=��a|���I�r?�,)L����H��`��=d�$H�'�ӌ�}����9/�X���
�mK�!V#d.��k��]a� D�|XxI�$��x�s���/��Ro�����4���Rݾ~�oF*p�L�B��&�=��ms -9�e
B�;�����~�,X�U;��������w-���~�������Μ*�ݶ��˦�7:y��*v9�ΊiVr���^�5Ɂu�j%쩋�HY�dE�Jjp5���3����Ú��~6��'���h�V� Я~�_6o�����mz0��'|�ɖ�P�oN�l�M����!�v�V� _�#@u��܈'�GAy�,Zo��a�2LyV\�'/��j��m��\�T,��p���u?�;(J���)?nJ�N�c�L�3�dA��y�R��&�]��'Z��(�q��)n��$x ����i��0��C
�!�D�+xWu�P^8�+�'K㲹>�	e8�BI/(��J�ι��)u��[��W�Ӝ����h�����Sj�8wt
B�SAe��@�����:��'Qc=�vz�%��Ue��G.�4%g��O<>_�ӗM�BR��'+6�Ά
l@�A��ƫO^c_<�/3��OD\ s��L-L}���R�~�R��Z�k_�ߺF B��������*E��ۍ���V�%xiz#+0�x�+��J�Ml�-(dHG�4���i�-ܿ�$�
O�:e�Y�I)9����7�v�uIW�k�J�L�peY�@�\�Gzy�t��$!y�T�����<�;��x���%����U�ny��94���ߋ,��4G����˕�8lb4��<�3�V�z�.n�����JX	�n�;��u6Ҋ�D��n�����dd�}����C��BQ�4��=OZ�Rب�_c|�fU����r�r�(��̦�|��>���R6�	[�1�����^1�<�Ȭ����V˻ٱL����T]yM�Ƶyu�1p%����S#�a�p}�5��1��u���EJy�=�����R�p�f��^��]���.��WJ����#��)���h�3̙AK�l<�toVeOK,R(7b$+W(}N�wg�ݾ�8���E�4(|E��\.gH+3#
_;��D��y;���V g_a�8�B~B�N!�)�=X�%=����@i�N>MZ�������j��X����x���������=^�X�����Mo�Jk�riE!�<�PDU8�nҜ\��z:�@�q����O�X]�Vq��ο/Ҩ+1��D�I�e��U������K
�Ν����Z\.�!��G�����x]��j#�jZ7��wO���+��">50dR�w2'(��r�EATw�{��.I�N����H�*��� �&�¨�)a�X�pEGx<�q����V�]���a��m�h�"�.7X[c%u�Ï<M:��5� 2�R+��B ��9�kq��n����]��E�rS&�1����t�
�q�}qq�Ә�2��3�"B������Q��u���c)^A��ֈ>�3ex��-�=�0����<I�h�·����ٛ'T�z�6�֟"a �>�]������=�G�^�r.�C�cيU3�a��OV�p��,iđ73�G}=��St=cP�(Ĺ�8���Cԏ���gv�w;������IxI3H7=!���JB˄r8~=w��Ohi)��ƓbT��/���I�e���;�����.#�����o�'���o(Gi�P7�O��e�Dq(i+ ټ@0x���}��>i�����Gk����Z�>B��i�� ɶQ��s�ׁ���D���QUuU'
�c��[U�5�&j�m,*-Rzr�6x_�������SR��-��I"'�Lf��owO�q�tS�=Hs�n��s����u�+�?
?'eB�W�t޲J��K@G}
1��p����Y$;��P(.���0_�hg��	>�y�[���A��~�ψ���[\|�W��]�+�k�5�K,G�/k
��rD,��������Pe�U�d2l�:ؠ@�#��-ً��EŁ�ݐ�$!�����a~�i�Zc�w�e���:5-g���s�����S��-�?r҄�'��d�o����jM��'�>�?y�/~��=�����j�V�_�-=���x�v)	�&�Pi�u�*���`XF��ID�`Gm-S�9ރ���u��Q*���e#Rc0Q�걌Gg�{��4V������$Ґ��n�"R��[�[�ꜥ�p�,����wznD=1e=��c���Ƅ�rN�}��!��!�&}0�	*�ϳ��Ui��
"�(��lH�{9�k�~���d=N־U��kn�tg)�Y)5�ț�4z����Ԭr˭���'M�Sk�>�w�"�)���U��VHUw+��,����^ͭ<����i��$O��R�3k��o�s��4>��˚�/�����&+��C�^wf�95gs-��w��;��	�]pl�{�MJ���u�a��P��]�L0�ޡ�һ�)��&�'��K��VX�V�&o�x�C\�՞O����Z=O&��?�h���tn!��-M�������.�Wuzb�+��GEXΩ9w���җ�:��n&X�VA�tC��T$R�(C��~�`�A�>��N��.��8}���\g�>4J�VB+@��
�bd�xÛFg:?]o�B���tX�- M��qn"� �o�[#��w@ue�
�	o�fZc� �j{�L�� H�s1�z����%�ۜ�B����-�TM�G�w��Di�pa�J��@��te�<!��;��}@3K{�~(�h@�$���5�wG&7m����=��8,R�WO*uy�?������U�ݭI���r�f�Y_�+f�Vd9���ǥ��J��㭄ns�_M+�������Tcg���aaYXB�N�`���������0R�(�a>�e��,p��A�P2{G�� WwiW�<��\vHLl��v����J��f|C���q�O��L�'#�;4�z�(��&���}�>	�5�����ckXB&�0�<5�7�L=�[����8�g�O�T{�A$�y���T�%VM�"��>�7���5����;��N��mp@�Ƙ/�?"�H��g5l|�량{���n�2�p>�*^K��=�a�,T�y		��z�:��t'������n%���F�Z�k�����t��ʏ��0�&�A��qO�n������~a5���q65�Y�R�	�V�gQnО?86��x�^D"9�PU"R.'N2��� ٔ��p+oB+�����O�o���
���_�eyA�ŗm���M���\�I#��?w,�D��ʍ�*IXEW���U q����牖@!H����7��Z����pǼO:�@뇂��� {�c84�љ�0�<r�Q)w1�U+^F�A����A��0p�0�c�(��cWONdm��Q�A3ɾn�T��Z}W��g�k�p��Ң���fL��ǐ�֑w�Y�L��BT�h��L]�,�|��@5m�/U�#5� kEfN�<īJ��h��by���
�`H8iq��ˎ�J+qQ#��k�m|�=��a�5��y0�D݈Z�è�A�N�jI��"�i�~�U�;�|��9���a����՚�m�Џ:k�k�J�y7?��n]�]�#n�`��-��S1���H�:�����o�0��s��|y�Cqv6Y�M�� (��CV���N��>Ҏ���B+}Rη�z�f�P&q�.���M@�Y�
z����Å�%�bPz��͑���N��a��5
b�E��̤6m�䝐i�q0\$v�_�bu"JF�H(�v>�U�np��S� �AW�?i�ڗ�kW6�2�ۜo:m(��dSN'����#�� � (�Ϟ�*�cV��!	���s�����q/csP2Xq��V�9�cYu����b|���J࣬c�`���tB��|먨�q�PfIt�6���(J��Y�7������������`�>�&#L2@g_>�=|�O�.�ʹ����}���N��ne:�~ݾ�I��&z��c�k��x�OK�f�������S�+;�~�ñ�:�X�%sS4�d�8�.��
Ջ�vn��*�_������p��>2�yNZ&�&������0�"m��a��zN}���
N�I\�BZK��xp��;GZfhy�:͓���p-6��riN%��{F �Υ��� @_�W��<��tQ�8��
��GH]'�l=|ؤE�X�ه�Ҧ�Tn�D.MP�u��wqWz�oڸ��9l:�x!u��:�S�gX�.`��W~��"���u+�.C
�/`�0�6�QÙ�}��j��j;�S����穧�Y�y�5�[���pF�u�=���A�R�p&8�R%��������l��Xߟ&"ӆz[w�Æ)��^��%�֓ɟ�g�Q�rg�����	h	���`
���P���+�?1�2�-�F��4�cY��[�F�w͍7*$~���a��;��>}Cۉ���o��?K(Q��Z�C�������o�FV=Q�f�77p+m�Gབ��41���y-x���_9FG~��̯>y�Z����*$I��L�H���[�ܽ!�{���/�Є�l,��<������?j��cOFG�S���"����g�`�8O�	J�~�z�Y�A����:%O,��mQ�	K	̀C�㦗1��|c߁�8?ՠ��u�|�)I�!]�rח��7k���2�XTݙ)#��1�EA��!@V���*	�;{ƻ�� �cM�>�,�L�zo&����I%3�M���&�Xj]�9�ຣN φ�� yq��8��<�"�f��Q\���͘�<+�@�" o�O3X�=���.��mH	�Z~�"��saUT�'���c�ܓl�NJ ӂ$��{�(
�_ ���p�y�BmU'?�zDX&q�+r�0�z�"3�Q����w�,f~Fg�H�����ƀ;�=��sM��NB3y_�*� VȢG�u*)����"�mF���(U�_*������$ȏԏ��U�'M���G��p~[�1B��9��[�z��(��^�N���&2��/��;Y��O��!n��V�K�<�����7�.��4}uٔ|G�QS���#�:��}&����J����{ m�6X�|3��A>���!��4�k��Yɧt ��N�'�<�Ʃ��-Sb3��x�&i>�q ��.>d�iI���TRf}��[�d��3�tR"BO���s6�M���=�8�ˍG�����s�1S�S�Sc�@t��p�Ma��{�ŋE��$�n����$����{���dLj�=pY@!�w�i('f5궪R��¶rz�EWZx׏�����(��V�d-�ޠ��O7�_{S�|`t-�%�|B���$���<���=�'z���a~Ţyd�eۇ�	��p2)l�~��:��s�m���;��ԑ,x&	�:����{&¤ɾ���
�B9e��y�C��ܵ����#�7��4U�>�n2cKdMR���V�.r܋�+[�Q�>�׭[�,
���I��R��paR�LʁN�.�P�?����=�f�V���f��(4�x?GW��J�H&#ju$�I��[�r��Ֆ�_o���ܨ��ͷfb{~���J3���gZ�=�y��#)a,9��ώ�]��.K�V�*@߳5�D���j��d�`�'&�ð���In'���C)2��9^�ġ������/vde;�
�QI���׌!L�E��1ؕ��sS�!5�LS������Ճ�Q��A�(��JW��9��Ha�n-i@Q�{.`���-��퓘nMK̵���OI"~L���R�l��s�_�{�p)�A�:a�B��K'<'c��'�L}����o��Q&��N�)@��8��.b`@M1�䉵�CB��~��<�U�{�VYU���U��q�]��7U�`���a.�몏pO?���C:�u�)~:���m���%���x�S��EH'v�y���
���@򍿒��N�n�uE7$�>���Q��Y� ���8"Hd�0�	�KY̘�"d�1+�\¾���<�S$�Y�&�L����X3�UԈ �ϟ��iGJ�Ќ!)#�Dv �>�����S�_%�`�8�ڀ_���Y8�% u��Ϣ�Q�_lOQ�Q�Z4�|�r.WtM�7C@��#�2q\hކH9v]�� �(+���,��99C�[B�򍴃v���[�Y�L?+��j��7��"w�f����Tc(s[���LV����C���n��=A���s0e��i��0ϋ1>�,_Tivw�o
�>�+�Y�J�	�auj� )��@XY������5��s7}�$ c�Q�E��y�� B~�׆�F!u��r�!���f�墇F)@�L��Qr�I�7��K�>3M=U���R��|� ��Rv��~�۲��̕���PU�'�u�V������s�Ho���`m  z����q	�?G�?�nM!��o�)w+�n�4\�R�����N2A�_AdD<fd8��R(�����{�ώ �B�hu�Ɣ'��p�w��h���`�.>?�m�s����$v���]�S��W푘�(z����n�'��<�ɝ'�gݫ=L|�xɃ\^
ܗQQ�9wJU֋�]e�S�wm���~�=�����z!Nhs�D��Qg?I��g��tI�xv���녾��z���B�Y��Ka`n�#�M��S�uZ��9(����S�����uXJ_�mЏ��Bg�/��u�+r�Y�rH"�����d�=� ��t7������zv2��&B�6|ʐx?� ��_e���;���t��ؾ���$=j�t��r�`M�<m!�i�sa�G��i��8X�L����+n�19ݥ�	���ʿ��8v�Q�J�J���h4r(ed��W��f�Y
�|O�ʷ:J � �^EyL_�|�y���e�im��e.�W�U���T�F<t(���Ѓ�M��f�;��>d�C�J�j�5�ZW�jBI�ְ� �54�C�l>>��5V�2~�4��M�oUf+���,��YX�:7�v�l�;�ͨ�B{ŋ��63�|��'���=�J!!9�I�7�F'������&�űP���_̜���D�?��H�P�<. ��>�G���F%P_47H���@]�AH�xE�!%������@�m�-�o!�$`���m3�*��~�M�5�j�O��T��3�̪���h	�ot}��?�1/��6p��٪]��צ֦�;o�u�X6��� pV	���j�����D����AF��$?��K|�x��ua��vN&���Kձ���E�w�qcR���U©n] �
�#7��3�㕵��V�jD�;�w�r�"�JnW��+SZ4��<�yy�)PoTnK��t�+�!z�ڷ�9u�z�ᵐ�R1���ؙ�a𼊞�����H�u�6N�؍�,WzЙ�t�Wa/���s_���o�%��(�Z�Vޚ2��Ԥ�04��Ҩ]�?�d׭\��nk�����n�}ܤ��l~��>j�d�5��C�8M�z��{[I�S�6�j��� `�d���ik4�8�:��è/v�L�8?�M��7�p����)�½�?��K�ܥJ`��V�2)�dD��:�P;�s�/W#� �I;e���8ǋSQ���}�o�AIT�Kؤ���Z����b�i+3�qn���̬T5;��i����PKxm 11��v�f��X��{�W]p������5>u��a����5K�*��nsb��8@���?.����LZ����|����<����X��p�#n��A3��F�Z�_6���XM��c�榦��[�U�C�i��y���ދ�DA�|�P��L�p��9�޹�V� !�#���Jݑ `�X�%\������Cw�J'7l�&��q����ۡ�?BÁ�W�hmV�
�b�yf}��?�Go���I��5l�l���^��^s3��������(k�hW�_�`=f��*Ͻ�3�&�ͳ3����f'�PG�L.�M��z��|X�4l�<�#� �Gu�C�
E]�V$���oO��`��%q7�Pb܁&+�Ť1�"nI����B���4�諬k�^y���Z{�����`/�,��%B�\I�a��\R����d�ҡ����_m4J���,Omp�%�������Gu����36Ԏ�H	 �=O���g\dht�V���O����
θ.��څ?��`�@����K�:ͦ�}���Pt>����Oi�Ss��5$Z�Fֶ`���Q{�\aeo5S�v�]o��"(�!���z��׆c1�&4���+ґ-JRu؇Tq��.B��ł������]�l��G^��g�K(�9�����ğ��I/�5]˺ݞ+���+~|w{�.���V/P
GS)Y)��sڧ��j�P"'5T�1�x�փc��Aˀ� �uR�������(+��x�ut��}<���`Uw�*d��֊�k2�	:����c����I��)/�{����n��SI�֚�Rj���R#����E�u�E,�����r���Q:�፰X)�����V��,ZU�s8,�0L!h��DVҵX�ٜ�9��QK낂.�������6'^1��-S�<�K�Wu���#4sY����V5Yb�h���5���>&}�*�f���>Jk䕹-�{$�g���|_��붬�k�(!�)Q�^�B�'Rϟ�]ɓ~�*�dv?A�wo�sU��c�jBtŴ���̝+���4
�o�cP�V+���<�����[���$��]�&^�sH��+HT�BZ�����Ưj'���ʶO"7BwB?�2�r]Ry�B�Gn���ܤ�O��i�O�(d�ǖ����@#�ߦ[W�y
������Zl쒉�i�K-��V飖f�fV��˦V��{"�̼O�G�J�#BwN{D����׍	��sS�#%b�&q~jl�ԛ�:�_��,O^�����^��eM嘯�����D�x]�T�4�>]�=�~N�9$���S ��W&󌻍�V�3r�[�^�?ý���q���(��Y.e_tm�`>�J�602EЍ3@E��T�Cq�;����O�? Pg�5�s$���T�Y�(��1�LO�w��ֵ�%@{�
�t�}��:���a�~e��K�T�[�ɜ��)�ӭ�X�z�>6�2=$Wd���+�2Dt%߶M�WɩnF��甫XkH�b�)�<B\�`U�@�`*��{�`���8�ί{^.�����o�
���?y%�pӢ�a�A��o˹�MJ��F�Uh�ì�n�b�+�v�SjH�8��\wf�0J��$�a�{��%u���hA����*p)p�E� �J"�uJ{(A�u�ڙė��`t$�|;��h~�7S��!Z�Y��ؔA6}X��:�^hQR�� ��W��沊��Z�i��جK��X3�d�ÿS
��
�w����P1��� � ��@�;5(#�_���������������v{ŝcBi��~��������e`�
��w�U�c�l��]��C�q�� Jg�rQ���#�3�!�{�f7�}��h9�ԩ����~	Ly�T
�zM1V]~�Q5?�� u�#ze����$�CSހI=�l�j���F�t�so�n�<08��i�%��u��=�Uz��9���G�׌<��8KE7�VoD^��'�Qk�h@x?��^�,���C=����r׽��>b\bWJ裈�r8�S��YD�fLoc�D,��~���<}�ܧ��k�f5�;���;�T�����7R�}�D E[�Ɓ
�փ20h
�Тvλ�{[�c�����S�ۊV�S������)�)�\ ��{�g���e/x�d�8�g^6�9`NP����L>R���*X���ƦG�5	A�c���
�B�4�S������~�2L&1�����t9�|&��r�O�:ۍ�+��F���WB)�4�9,�E�z̈́Q�(��j���� ��)� K{y�
qѯ�\�P�%@�4��ͣ�	��˕G#�I)K���m��S憚�bz����d���Sz���U�M��Ȭ��>#��^�� ō���7���tY��,��xth��si�O�dz>uC+l�.ݩ�4V��O�g��E���s�B����@J���<�-M.;�^t	����U�#�=x3a��Z���/���{$�%��5{�`x��ѥǄ4�[k����n��w>b�,³�#�d1��_��1(׃��Co�!COD��
@���7�.�Y����Y�T(3�c]1C*�Ȓ�������f�pxx��s��������7��V�ѽ%7Uݴ�i�(�;�40-2���Љ����h�uӥm���\W�4�p��Qm�P�\^��E��������8ul�i
+�����y�X7��Xn����w��b������@��L��X7�(D��~]�+8�3a
C��¢��.�;w0S�р��8����z/K�,��.�ȊN�{�!V=L�`Ë��<U>y��"C2�o�JsZԀ���]?�S�(�Ԥ��*q�C��oJ�: ,R7=�j	����2�$sw~Sb���ͳAʦ�����8��{����&
G���P��&X�`�+�ֈ��x��3�����Ny%�y$B���N�<s��Go�4~]]�)�D }����������yi)߯,n��@=_�)�Ml!{8�X-�����m:9�����v��Φm�c.�����fp���B|�����6k�M?�i�J�X��(6�rE���ȓAL7jo.��<�f���L�.B_�(���������9;Ay�{2F��V�����hK!I&�(Q9�����!	�`ll;��+2�^L={�j8��=Ӧ0�������V�K ~����(��O�j#ߥa��ゆ9N���h��s��f�3��(�\l:�olP΁͍�$rE��:�"���B��vfH�ѳt�:\��t.���Uz�������kt]�hB��GE��%qk
���%�U�ΔR���Q`0�2:<9k�����|�28��ZJ��O�q�ŉ���腻ڢ
��a�����UԄ�E�ǈ�G��
U�w���8o���p��b��T����:�.��0f��_sq�)j�1\kh
��i:}���9�ZsHz��)��qvS�xM�%2r����5aw�w[��6�C)�-�I4��w|d2b�"����0�����Xܬ���G'KA�q�~��j�3���pX+,�v-t]\k�!G�Pf��p�,�u@gEu2��?��n�I�l�C8O���e���CL�[)r�8Dt^X�<��p$�]��jk3� ��3�wņlj�_�O�І�\�2]�x*B�C����<��mP���s�f��A��k�*���:�q/"�?��S"�*1f�����Q��7�چV��@��lD��	pơ�ߚ�{������|Ŗ;T�/p/9v�Ɉ�ɤ��q�z�3�j�����i��&g��z�R/� y� ��+���.E���}���G\���:���f�Ι���JO��a���Hƌw6���|���|����>]��.ؔx|�dRc@%�n<�����=���$�x�=h,J�z�	�3��|M�IE#�2�U��Z6�B[⠳�Fk`�B�|ú�%>u�S�"1�P�Ky޺�ˡ6��!��m�J"�>��U��ۄ����#c�@�&��t��J��^�����������e�g��n�(�_���l8?,�UX`~:��Zy�
���֮���l���DP�L%e�d�Q��d��P�p�������'E�Z��0d_S��_��W/�k���D�`�'���{`��U�H��J_k���ZI�����#4s\;�0�qY������� d8l����>(��E�
��kV��@����~к>��}��W��M�7q^`$���� f���G� ��2��,��=)��b�����C6��ÃA}y�4��:H�U�>��w\��ꛘ�'%ăĘZ�9���p��m?w*s��ӣǝ�� B��F���J�)t�_'2������r��Uy�}�a�x�:�b?"����)���L<w}�1�q��}��@t5��^|-\��h2���t�8mpsnS�$����/������$�"9Ds�E>��ެn��^s-�J�#�����]�� `�wvtt���=���ҵ�y)�� CV)��,��nLhpI�JAɤ��R�vn�h����J�Ν@��pR:�\����+����~C�>�<�\/왩9��M���$P���l�@��p�D`.i`�qNK�3x��n��[�D�5��9ZQ�OX���p.�䲈�@ȇ�+]������l�O,������i��e�Y���@�53�\4�6��ed�e���賅i���V�)��X8���1-���$ qbsŜ0��'d<͈�[�^�;)��2���}b��yi�O �y�m�{�n�r˧���
������##���R����^q4����3<��m�G��'���"'RQRTXW
#"ZWؿ�9���� *��#��<��g�G�Bﬆ9�:ߨ���x��0�� rvMj���W (܍7H��K�$y��vkw-�?ѵ8f�F�Hꊔ�<��ѥ��}@aO�A�����hZ�[�L�Xt.�q}0z�Ҹ���[6Q�p��I���aP.3.35?)�nk�k�@o�m�5�H}���ܒe�a��Us�Ȫ��7X�a��k_�6��@f�j ιZ�<zY�m��R[,�y���+q�	x5����5 �1r�Q�)F���%on�gA8)�4�\KY�)6S��}��ӑW�Q�u�\4$��ډ���r}���j^k�-$s��.��@V/�x�~��@/ )�پQ<�v|�v���|[����a�y(������S?k~[�}��{my�9@�լc-��A�߭M����-�߳�����zH�d�Y�uL�' )�'�gc��@��q5�粄EX�9��3���i͇)D�!���X��_��Ek�W��#�^�I�G8&*kͪg>��QL�K�f~r�숍�j<���	9�(*A=J��{w�o�T�A��Ad���q����zT��y�6��Ƨ*�O�/��S}��Ѵ�����h��p�/pU�~���/��O���ZRA��
���[���ܜg ��p1�J_��JRpra�����=5�:��V��>�TٕޒS��W�ztqO) ��@�1��N��k.@��i��1z9�7��aS�u�J���:�go����u��~����
�D�$��M�_�^q�S�!��.�Q@t�� 
5� �։��H����(� ?���*u��f�ޏ�E+��ky��$i]#��K�¸������[p���o��s6غ��u�N|�%�>��?<�M�|K	�xt�,Ѡ~_q�ݵ0`���P/�l"T�����w��+��R�Gib���^mz+�񦙈�5	]+m�F���x3�ӝ���������v�I�Į���0_tN�yǪA���8?������îy;ǜo�$+�`�:���aS��p���^��V,���Ew��O�l��@�/`׻g��sr@��/�/T�vO��ʤ%��n�D'\*�Sɮ�vR����9bu���F��Uw�Y�Ԯ���r�˖�z�0��	�(604^$U�Q�xp������Xb��a��%��h�mő�����V�X#�#�Ɗ��y�[��3Mw*lt_?�Qjz��b	�"��1�/��	:���Q�@�8J�H����:DQĒL�=XQ�^`�n͉�#���e��H�'�ӾZp�<�Mdnq����b�;�˂;u^�bXA���S󯥫W�j��HT,K~cUb��[�}���D(��<�.WRў&��F���q�x�i�.�Дr+�߉	fj�jf�?�����
����D�2�'�iC'E!|ȸ�� @�6�mEJe&���;J�W�D�/(�YAG7~E�;���!݌�MbRK��M��B��-�	����;?J��fI;�-j��+��o!�,F
h�����_���M�>�VP;�m�O��Ơ�/i8�Í%���A�>WG�	��6~`�1�f]�V/��?�Co1K��G82����=�?�?m��/A�BzL���@7�m����sG�ڟ �.��vǉ�o�
_���:�+T�Gq��\SCku�4�E0��,����=�e�;C�r�`���To�P'� �9<�u�&�k�������Kx�#+BrB�M2bt��0�w��ǣ�K3h�������4�\m_��#vA�rV��q��6G1i���龼�鬭�cA�+e�B���������Q�&\+eq]��z����#&�b6��K��󿛮�v|�&� ���&���B�=�,�>�ă}o�&E�鮽�֧�V}�"I�2U���y�`��ٸ�K���6f5'Fa9�!;�p��5Y�qz���Nh�z:+���"��}J�!�Of��\w	���p�P27N /`JR5�NxD���H�
j����\����T�����W��d�����!��}s�1�S%�FA	7bC)�Dܠa�[$}%(�],�f��$pm"Ɛ��X�h�-�!z�3`YF�c�\dgL�LC����e������Z�+3������O��� QΝU��Wmύ�"�3b0�\£T#�탭�����ݰ`G9��|�J�	
�/���� IRt��U��u���@FZ`6�lS�$ج�w�Nw!	K�w�;�����X��d�С�Q^��Ux����?{M��r��9��2-�e�F��`��pꆦ,-�'	*zT܏�p#��d�iw�KW�������Srr���FLJ������֛껚�luɧ.�o�%��L�^���]7������oՓmb&�m��p�O��w����Nh�&,�����dT�����x��>-S�|h��K�<	��Mm��f�k�̽�~�8	�	Z'dVL��in��E�D~���mO�*��cb�s"���D�X͔�ϸm,���D�c���L�;�=�~�uy�ȏ�,�Cw5����3�r��gd=����.'�BL<�s�LOy2�	E9[ts[�-/���'z��	�Zm �"(ۀW��)w?$��"��QV�$����H�I��q֮���р���.�
Y�I��:`�%Q����Q��ݧ�~g>�_���w�X�����g��I�+�Fvσ23��]������%��s�N�VnOO?���ӶI����l��rz}�\\���F_=B�l?'3���?���A\���֐�i�MNi�n��f�Nu����,o��>�{R�S0		����t����mU�l��2F�46�f�I��"��t A?_�Ab'�6��0㺡� 'Mb��c*c����I���B��WF�E��$^���d���6��Å*9�t:��uY�����W@}d�"��$6d.LZ��O�e����Αr �=x�Z-�tǙ4��䤇dcϿ�M&R^)K8q�� tl�-�����>�O��X\P�5�������[�0���*�$X��pzܠ7%�=7֯�sy�,�T��[ӏ�c�trZ\���-���� 8���a����Bt�<P����t!�~�8��`�}G��ˀ�Ң9��y��ft���Wƙ �ԗ�:�+��(�c|��a�?�y��6��Q����\-�g��~��$���7�TodG��X~8{֐X-~�D��?��[�z�"�
�u�zi���QN����c��S��LW=#s���I�Q�:��,���l�,O���&�Q�����>��3���X�����.�c�,h�!L�C�0K�-x���]A��6
���Y���	3:�*+h�R�$WUbJ�i:������
*$��*����N��T'u�5���:EZ]$*Qb%���W7�z��ɉ�L���
��>I��A�W �3�w|]s��ڥa�|�G؂���|[�@^�c�@�mr�� �Tl�?��hqT�S���֨��.*�~�Wj����Ђ`_+�S�-� -,�HbefH/A�`�z�O�B�ʚ��"�0�<q�^���E�� ��47��r��1��#��ک���;�w@y�`����V'��u)�$_hΏM��X�O��њR������]G���켣4I�"��+W�UxN�鯭�r7E�s��c<��y��8=��h!������ǡ²���I�����
�exJ�����3 �0�ҕ���:���㈡��.	�	���&A
����H\�@�P�v1�tu,��f�/�����Hﴮ�V]K�.��d��k�X�CU:��-�
�\��.PL���]���K��[#B���)�i�̶{B;ZM�DA�,j���I�xf�n��lަ���Ó����(�l2�$i�Uy���.����	c�o2���i�O�wC�l��0g�����\��N�꬗���
cY~>`�Cl\mn�=OA��)�c��=�b�O|���&�Q+�8A��ep�:��W���}n	��T�41���/ь�hraj�e�wj�Fs�8�4�.�ˏ0����	N��)C�zFd�E5�w��ZB�x���Md4�>���ٿa�J�6�`#o\_IP։d_9�2/�hzB�F�f��B"z(-c�y���h?Aiu(�urc�ὢ�5)#q�\hi��j�^�|�#�����i!ګ�bǽБ`��.�t$=	��E]i�/;a�q$�[U~@ɫW]`ej�!�f�ԭ���-[��_w9�d��1ij�2��w����?��&=��d�٫א�O����*�E�I?��f#�in_���#>��<wo��
8�>|�>Nʺݢ������F�M���5xh��G�W �@�7��G��_��X%w�>�XU��-�M��L�-�=X
°��l>�qE��n��vZ#e�ה���kj1�bD쟒�`�:+%f�E�����K�Dy|d��A��>��� ��y�;Qz1?���������>������m��(}��,���}ynA �@I	G�z}� '^�I�Zm)K��׈����|k�(�R:%,4�frZ�t`�p�jN�{IzJ��
&��B<�op
�a���]�L,� �>&���� ������7I��q\�#O@�[s�����P*sUI�$��?/�����ю�g<��x�Ryu>�M7_��ù��4�A�%�Kt%�Oq4xϣ�����|?��dqj� �˖�e9D_����H�zjQ��c�,����7a��(��CV���O��I��������~H��ٿ�P�z�M#h��.�]�Z�N��䯐�.��'�bhoβQW�YO��=01L�>p�э�p��<�S�4�#��H ���lRt+��b���i����	w��}���~���A�5��/��W`���@v�c�H<i�T/�A#�$ļh�V�}����6�&r�G.F������mB��*�P��,���qүͭ�i��G �(�if�����`	��݂��L���9�DF1�<�.vz��-�B��`v
��z�oFC@u��R}~��P��H�'3A0��V����2�Q�R���o-I;(�U$��t�su�<ؙ�ĩ2�V\��F��(�Ji�s�B�&��d���0�ق��iQ��7d�����D[?��n���PA�>B�bS�!�Ps^h1Ҍ�����{l���������&=��Gy���g�)T�q~2N�[���|�L��G��Z �"]��Ŧ���o6���_�V�'�ڔ�h����6�.�
�>�h0�XXs�G��De�B�>����C&=E�x�g��%�t�����M�}��HN�`k$�s_{��K�WW��������ߦX���1�M`��)�%�)E��R�APX�Օ����/�@ )a�5ig�R��5���VɄ��x�H`w�h���idL��9�N��|��VU�j��XGl�H��[		$��>}��#nj��0p7C��oZ�F����h]p
8�c*�l;8�e):H}Q���'�0��!��J�pD��A͍�RE#N�t�;�ȕk����XK��(�������r�
�;��e!O� �[qp��tyi%=ݕK	8��^^�Ҁ����#k&�_<�7�Џl^^f>��^񹼉�(�L���K�c�cн ��#o�w�����fe�7Re@�8�WY=�G�¬_�cß��/�`]�P�&�sޱ�u�$�%	�w�J��o2�}�d����Sh�!F�`�m<��̝�U�����M����;��c�7����(�����Z���'��Z̛.-u�zn �s�k���m��R��O����n���=g�x�5��B�n�G(�[�a��X\� �@�E;x�3�_½����؎������hty_|�mtS���t���&���aE�Ӏ�G�e�ئv�vo|�OᏫc�f����QXzi�tU�����/}��l��ѿj��y�ꕤ��=�C����:�@P�'Õ�\(��D�(�s$��@}H��)��M��۳�����Y�2r�d����k_�����03:��O-���M�V���<"��쬫��q#�Jw��N�@��̡���Cvcܰ�݁�$z�^�6mu�\����80�	�qZa(k?w�y�W���¾��L9�[ƠI�T�<N�\j�$oN��m8�ɔ�J��U�깢O��d X��m�r�7y�S9:�͝ϩ2�&H��\�|�ոQ��Z6뮟�u��eb��� .�g"�+W38}b\�s�oQ0�����8#@2�U�PT��P�v�x8�WJ�FP��	�X��Xe�o�XI���5��MD�̉S�W@b'e��黎�!�4~wu��c���u��]ۮ���_�.F	W������,K�4A±|X8�5QG\�o�K��O{�vn�Q=�%������!����I��n
�׭��om�����=y�Vǻ��~�樶�}�c�-�FiN�������)u�a�O�5qWz����6k����N@�	񰭌�z�a�`j`by���I��0�3����Ƃ5��(��|���,�y�����⶜��ɑ����L�
Uhk4��*��yɘ���R<X��,�Q���\HN��o�u��ڥQ~���.^ຑRb�#'�˪��KX��f�z/u�ZAA�`O$c:��ds��	˜|�)����	��M������/����;�S��z�(�YC##��o�3$
nP#�u�Q���;BM�L������=>�g�f%W_6��2.��; ��"���W�(cP���2`OM���vn1+��b����6�|J���~��߷�x�Xms%/+�/.V�z5��ӳ!���.�� �ߎ��5ז���]��&��$��7���
�;W�� m��Su�r�*�:ͽR��H1���|�����L�߃���=��ޏa�͘Znfҋ�sAA�B= n؉�j٭	G�ro�T+��oTꋿ�į��Zs����Z(;���)Č�"�V�B��~+h�̠�� 0��DB��j�I�N~�� ��
�ӆ��(�"K�����n�au�� k�)�g��!���Q9�w6��Y�I0I���wĞ=ZTa��5�dM�A%X8��u�&Ht�l��-���[�fA�����w�t�<61�� ��&߅#Y
��o)�s��A`R��I�>�|�Y�+t� V]*%q��(�i�ki����T(�[�=���Xdr%���^	����g���l�ӳd��$�B�IbY|7{t�;���`�y�-��˺�*Z�^b1��v���Yc��P��_vک_.��h/(��8F֠���� IZ_��OH\!���5e�,1��:$�B/�A���R���@����O����;}/�*��LX��:�����0���՘;���)�n��D"B �,	����]Mm o~�-��@a��C�����.�z�/$@����'�e�uY�P�Z"$1�e��^Pa����.h?K�4|^��%�`>�Ւ���oA+˛�Š�W�Ou�����$�D��ڞ�� �0��������Y���L�-x�a<��I��[\)�
=??�>����'��u��}#g��&j<��zf��mzV���2��$�$�f�N�a�u�F�M�3�>�����������+�N:%�����]F�������q!�H6�/��h)���S�pm��r��{'�|�^M-�{�4��9x9F ��U\������i��#�t	 ����	_Xs�[�9����N]|
��r������(�M�y�(���o�/L�Ҕ�l�ԅ� �喀&����&+����M��H]&¹Dh���'2_&�����`�ҁ	��R�K�(���US4�To3�:I��]v��q^ʴ�q�@�!���ޛ!�-z��?"c0ah��W_qLς)ɛh�����)�#c}zRζL�4f��������E���~[=�������E��V�ǣ��/��E�A����$>U��a��?�QzU����Թ��Q��@B���+��KGh���ᴉ	U�(��tᡭ�WB����O�w�=5�5��2V�ƀT��"�1��$�c["��Z9��fVp����HE]�P��]���t �ջO#D�(�(r��f1�9�"-��ߋy��V�#�G����b&Hj�wX;�R�O�Jت�&yry8`%��Y��M\�)���O���Y3����8H�R�O�o�~����g����]���ͽ��he��m�v�Ґv�n,�R\�4��i*���?�t���i<m6�D��;���Mn>@Vy������-���Y��s��1�!�Y�͎�^�  ��If���^�w_tP�װw�>���xw���Kj<a�㕨��!�ʗw�b~�@)���ѵ���E'�]}r� ��'�}zt��t�(r�U�/�ٮI����vx�@L�+;����:��}�F��
w�҈����}OE�����͖�'m�hX�(��<9U	=�`�d5�˾1�cN�����:V�[o���+Uwi��e�vE���t�ϜBm�i�m,�U���������u5UBUY�əа1^:���4�(BO6�K��B%�����6�Υ���_ͣ�����?UO�׼|��s(�,5̓�E��M�O��A��[�8D����!��}���6�찣�C�a���M�wT=���gw��@'�Ժ��ѤW�]�!M��:�%�_�������v9�7Q?�ہE���wpu�6c�5T����V��^����4��HZ�� �x�N��E�*�x����4܏��|LŶ0;Kd��| �A����1O��2Z���0#��n�Gay:W�5�ZK��a_�p���C���D	 \�E�"L�0=�1:bbX���Иso�9���ǣ���,���>�F�1��Y�&��^GcM�5�*����>�|M }B�w%v������u)~��G�~�H8��Ez�\q�!��5�;(@,�Og���2��C��� ���!��C>�(�Ů�͟W��#�p���T��ߛ�rnf64_A�	�~D)/F�3��2~�n1�尽of".��},-�:T�A�H�-�$8�~��}�EO��p���&��pG�,�����W��fA��No	���C�=�b�!tC�EmS��"ߌc��e�φ�45f�>4t�t��,!P�}"���F|,"<���h]�Ƴ�����r���1@�trr`=M׮"����X
1p�\.^���v8�I�jn�/.���v���7���u�se�+���͂ŉ�7%{�hE0�S�GԀS G����\gHR���h��:�̠��l�V���Z�5V`�RH�q���Y(JOB(F�ʫrS���U����������
L?���sS�{+������;!	��_	a��kE��C7�]h�c����`��ў�,"��)aV*��-�����^��@�`W��҈ܩp�@��=c��ciȌ�q6�C�0X�CZ�F�xN��.VCz��j7=�p֑ro�	J��'C@s�0�җ|i�3G�`{�/���@XƮO ��1�
���\�ؑ���cN�	����^K<��6/���{)�2>2�"B�g�b�Y�% �Jf��!r���4�h;�ZE͛�r��62��כ�����)���w��Cvכ=���8D�zycK��������-�������Z���aB��4f�����)}+P�Dܛ�5�M8�G�rOr8|y�U�E���ve�0<�RT���B5;!����k䅞�[67G����G������s��xw5���[�/�p��V�H4��T��\�Cl����Y����4������BU緤t�թw�w��q�T�:��N� ��kT�w{��E~l+7)���3]��G!��V�;-hc�j1����|<�l���KR���тiK���t��|]���'^uXp�zEp���h��r[qqv./e�z�n`]�û��$i0yaٴ-�5�`�fj�6�ze\\�=k.��b'ˌ�
�r�aCR�e��;�������蟽�!���1�,zN�Ǟ���+������o"��3}U���������K����&I�?A3@��`�r��R�ͲH��X�ɯg��+WN�a�>j��MuKw��-��G�>���+��3�q��ݝ�y�{�83��0y�W#��ո��=s`�>Y�J�}DS��׻
-�>	{�������V\rǛ�2b�m�\;�ڴK������:�� $����T\��b���Ax�w��9��u� ���lM���ɝ�y����d����0"r#�n9����������h�e����kh*�Y9@�]/�o�xdV���6��Ryd��*��OfUx��Y�I5=��z��Q�7&U}&>��5�i�Y�;�!o�a��0Q��WV��?�e=\r��W)+�ԯ���3"���_Z���,��7�i�nv� l�p懀<�Վ�U2ևj>\D�y��z��mx��q�'Q
ܥ��:X�h�	��ĭ:§$�%����G��=#�#+4�`�9�~�,���Lh�a��w����iq��1�Vf��N֑�����_	���.ME&��4�+���|ۻ���k�3�u[��=���M��}��Ɩ�q�ߙW�Й�Egr���H�i2��l�@2�ۇ�w,�Є|�̜��T��p�MX��c��B2;Ҿ��_-�����m�u���[�� �䖞� ����[�>�1�[�u��)��K��/h�����i$�vTl�^.UhF�:�#9�J��Ny�q���5��4�gӹ�(���Li�ȩ���Ӣ�ph�����+����2�.P���?0���Ӱ�i޾���F����^��c�B���(��v�{�!��%�r������VPlP@�]�^�`���9�ij�ȑ��P҈
��vCU��B@Jx���Js�6��0�kp}�@���A�N�8�?����V��yR�w0�L؛�JTWY\L�w�˖4q��\�Q����s!$���T��������}�%�2�+���V����y�1�u�DLP���y��?2��D�S^jg!�/_(<��(��)J|1�s�� ~`>*�E�F��BL�#�߭�<�5�k��$���6���F��8|��i1`�֛I�������Dy#JAZ_�G��q��iCq[j����&*
R�J#Z]m�q���m��:�ɨo�uO�Rfֺu��۬~��d�5X6h1ۮ�$�4��w+�V(� �m}����Z�ѻ-�����(f��O}�]�����r�7�������3O��@�[���KO��n ��-�F�',��4',�I?�Z���Bw�]	�*�Pjs)���h��.�}{�'�V1莦���:�˵/�N�ԝ�G��t�3�]�k����٢lY[j�V��hL��䰵���YE5x��x/���8H0�fU��y���-l
݆n�]�ʾ�����p����껫s�c%JS,Uľ�)u
�]&A��I�����
,oN �E�vb�����Vy%D����qW�9�:�<�l�fO�<z.oTa�R�nb���� f�ci�3�q��ȯ�r>�ݜ�%�������$�?��F���n�>߫,���c�X+ݚ����{�3��j��*��Ճ���ƥM3��gS�R���:��څv�ꊇ��i
v5Z�8N:�fL�6�7�V� <�Q|�d���V�;���ТShRdQ��4M��D�bwe�w�T�r�*ٲ#��r8f
	:5�I�K�
 UU'#8��M/+�� `��3<��!f�Zm�B�MS���iӒ`��Iƞ�F�|�)6�'�8��:�_��;��47�u1�q��߸w"\eЍ:�a���gG7t��#���Sۃ�-j��/��:�g2,å�&�b��s�LN���x���WW�TUn���P��;�6E�F�Ԁ���K�\�i�F�m��HJ˛ΒVV{���KL��B���Z/�kL~�� ʆU�td�]�g�8�/]�m����P�Q��s��ZY$+{��<P��+
�w���<.�J�h���YI=N�����d��h�y�E(��>1uF
Yt�ܯ~��'
O^"|Zu��su�`���F��2�������1zԨU�p�y�ئW�-��"�y�lI�Qʙ������7�C��h#��n���-�̆�O��>� �p
�\�l&{�?����"62�K�]�Lb��Tv]OP7�`O��R��߂�\� ǡ�s��$!�"9ͧ���j�<0Q�NPs)ܷ������%�7h\�b�-�T��,Ѳ����Q�9����h��M'��Z%H��f#+�9��&��6�,|�Wf���5ǚ!������;�^�>�_O�f�~�D�4}�,p��Ul�.�^!���;�/��D�L�Y�"�IA"VE_7�ѓ�Z<<1���m�M�B������}6n1���u�Ht���cJm�M"�����J�
s�,t:�	��G������	aO$�d�9ǯ:W���'q\�3�
�嶂����0Nց~oUpZ�H�:
@��C��5��/a��jA0�e��Q'���sv���M#���������p/�Rx_XɁMK	9Ԓf�u���A	|�/��Ü��k��(�I�>�i�Ny�)�	Tm4Pt��I�'t2�]�a�A
�k]�ܹdm�=����͊���2+R��v3��B��!m�������hr�)����M��w��v|�_$�ѮWC��j�ou���S��>^,�.
D����F�z��q��������?%���rW\L�^�:�y0�y��X��V�#A!kOB`ס K�y��+��?��8T�T�/�<�c�Q������Gr8nL{t�D_�¤�l<Z�L�7Əl���m����Ex]�}���<a��˸�@�q�D��ɡ2�m@�Ύ/�է��1qaF���N� �k�~�$Y|�+�F�=�p]I��H@6�of"Ǆs��P�=^)�����1K���Z������&����j�j�lZ�ǆctR�׊����Nm��*��cF~�,�Y�2�o~d��7��V��q��ׂ�]�lOɘc�hO�?e�~���
��>�)W���4̗��� ^�n�>PX���I&�#��'	���-b.{Z����5��B�4K���� (�2'����]�� '�������3��?	� C����}(2����u�J ��!�0��I.�^�(���A�P��}F�D�b�~����g���
�f��y'���ГA�!�=G�de.�Nہ��5ۤO�e�k� #�1Tq�jF��n����\����j�"���W�ڟ���߷��֣StL�_m��9���_�0n׃����T0�1mI�B_�!mg�a� ��(>4>�lv�SA>�=׶��w������j~K���\t#�P�\. ���ͯ�(��l�hT�$)���(�R�ɗ��q~y�a[~�{@�`i`�y� 5���m�a��M$q���xS���d|'o��aT�E��جki#���Ļ[L	�Τ�3,g��(vO�p�a�`���[������)�^� ��<��7+�f�&O�1:����y衠�k�G0�0�ţ����I�ԍ�p�+g�dk�s�93Z��WH�2ãx��X���IKr�.R�v���X��D��67`,�F��5�����B��B�'�j]oߴ4%�AI�j�W�)Q�V~����řt��n2 #�jj�1�0KT�%��̕��S��+���l�	�c���
���3r
�@��f���{�@T��U��h\�d�v��D�����oh�}h�Dg��"�>�%ˉ�|�mҲ�JX�\���h	���aBB�@���%���zSy׮�oV�[	�`�ܣ ��^�`���;��*���]e	� ��ָX��6BO�W&u�)��']5�u8KPm����g�G���bЧV(��B�`��`����+��~������?�{vGJ�[O�*���I��1_����Lh��+L�Y?��!u�5Ld�|qcj+3 h����~��T����O6m0����H.&�:�T�v����bO�q�:����xݡ�h\ɓľ��]]��:co;�	;�s����4�p�&�t�N��]6��7�Q� �M�B�ȼ�(P��˒�1 ��L�H�Ψ1��v�P�q�Dr��x5�Y��#��lrx`ju�-����6�6Ƈ@���2Sl�9 �fy�9��M����2v���r�[&S�P��d�#��lTJ^��:̠���;���?ض �9yVn���9�=[:���>�w�нi@ht�Hm%p��7Xw�2�Tq�B:n�~`��|�b�kj�8�@=�&Z�V����������}�ۗ?Ԇ��p������@Px���|����3�n�� G1m�K�q�>����gv��Y ���Dg[�1/8��䦆�zG>���󳓈�����-dE��(I�|��n�T.�[,r�|d,�混�& q�E�ݪ�!��M��%ۨ�Lbd����W��*�8��XՠI5'쭰�2�rs��u���7���gt7�xb�\�e���i5-���>2�qŲS�$;��w�'����=��5@�jR��ݐ�J�M*���7���{8G8���;Z���=ԁ�̙�������uJ-<Uk��v2�� �s<��N��|p#PK �`����#N�����|��p @z0%�g[Yゝ�w%�X��Pqa,�����X�2�U��P��w� �a�X���u�o��"J�C��i�[�`t�=bw��V�.<�c=m$�)]�㌣W��g�C��Z�Rc��!����rP�'U�}�ub
�k #��e������ãT܏H`���x������>��:�0�pp��p�&�tuϖ�`�\��Kg�(��{Z��+�c^�`�M�&$��*u�\aN'�t��I����l��"iNJ�ԃ�Ҧ�������OxS��Ʌ%�&��Br��:M"���u���a��.��Y��=�<л��6Dq�w��&�~�����`�4�"��Pu�.�y�e���s9�-Ǻ.���t�_���G5Ҝ2AF�����v �(m����v��2�F,�1:x�ҿ���<Y+�^��+��FDooP9�+=GM��LI�Nӆ���@$䳂��5ԛ�ک���
�>��vښ ľ�^�@���]�]h��?���V46��|%�����|�r�$f���
Y^Y���]A�媲�PY���CK_H��#�v7�bGc
oX]ÄZP�w7�\�?�A��~Y�"���]�9=�*1�� Dg,��M�˯3���lE^�Q��V$�C�7�wQ���}~�4�.f�Ԏ_-eC���	�,4��e�y�y���c��Y����5�)�]$!��R�/����Q��V7�z���C�<�Qw�]P�B�VW8Դ\5����'c�h���oJ��|�o@F~�(�X����=��a�bN��O�Ŏ����ٗ���@7#�5���͏mR^}�t�ћ<�I�Q�S�C�Q>Դ?�)��s��$��@�<ke��M/��6D�B�_����kF$��f�$M+�[S�ĴC��.������������jj�1m�FbH��/eg��[�u����GV�c�Q(��8,;�?�Z��\��&�`s���g�G���p7�������U9D;K�h	�;��f.�.��9��Hօ{:B"�6�v�S����OǰgR�3#��ToH�.�rġ��{�B��Ӂ��l�K�9��&�Ul,6��-_���j'WD���߁��λ�$c,c4}Kv�V��`ݗ�{
�U�Q��v�;9�=2fV�jL�A�t˾Ǜ������c���y0�|?���e�I��r�x���4ZM�U>�Y�E���j���E��fl��*/�FWJ�ۗ���ZE��yn���⺆)oq' �y�䆈p��i�ߏ�Õ�_IY�1u��\Π�<��	TE���u�,�B
�`�ȷ�ZJe�M�A�������̗,,�(�����W�0��v��K<A��P���ot�"}Ξ�)�Dc��6]6���+<Z�[��ਉ���cڂ��n�
aG�Q�qSK�;���)�~��7,']�Aq-�w(�%�s�cn��� �b�z��EہW�,��nED8��)t��`X'B��Nk�(��͂��ٺ[�:+x��ſ1~'��s�w-$c��#r�t���Mt�!Ǽ.�؈qt��M�P��zﶁ���pp��>~g�S_$9���f�C������U��+�[�\��i'�cv%1���@�없������Oʴ�����w�E�^v���`r��e��bK�����U��ӧ��c"��Ѽ�+i�2��~@��
�ۆ1�o`�loФ�G������l�J�|��	�=��>,��90#�3غ�����L֕�'�p�X��\�Q��1���tw��1z#ޮ��ؠi�D��F
Y�]��,�4E���� RD�������U��5����� �.�9u�L"[~Z����Ę^
���t6�u�\��v��	3������D�������h�E���9�f����ߡ>���Ь�w�Ѡ�{|!��HX�+��I�������F@Oܾ�O��"�75\J��ĺ���U�;��8��$���0i��A�b�&l�8��eq�Q���ߺ�9ql�`Rge|�_���D�p���&��"������w��XO�nfք�.�`0����Ej��-Ū}�]M=̓��.�����.>6~H4��+?�ᚵ���~��T�鿘"=�g�V9%�<%p�1�AV�����頕6�M �2�V���W���(�@ǝe�2�~N!�(��A�+����H렒��nSd�w"%Dק`
����-fyz�f5�˗Z�^Ol�&e�hP/��sRc5� �_��KW,Z���l��h��h�ؖ�G��Ҽ>�A$�Z�����F����� �mQ#�g��J�حJ�W�����o�G,��H%SD�"�By���T����ST/jK�H5<،�`)m�ѿ�?'Qeǭ�hPϯT��^Vc1%,I{(q$͟��Q��3��&����ǂm��)8��x(�h���p�4�D�ˑk����ޝ��l*�EHͬ�X��r%7V[[���a;�RgiA�l!�x�Qa�`w �i��\\8b!�QD���zUVE����ྠ�'�A�P]��$I v�l魪��r���W1�,�9�lM7 ����r���7���=ޏ:K_N �д_��q�bg~Fk���
�����lID��#�j������S���2Ŗ�����1��K&�3�E%�B�m��4��f�Lk�D�=��"��#���>������i��묑QhDdY����d^u���������HT�kAA���J��>Peت:��,.u۳������(���g��U|���)�i�qc���Ke�禑�Қ2n���՞ȃ8o�dvYz�vr~q:*�{�HUQ�N�NSP7�>-��lN%�8��Na�Cbzٻi�w@�[���c�:V{��U��f�KZ�"gA6�%>�x2�+�����ͫ ,w��)�I�_c�L����I��(�)��,P�"�v/gTb2C��'WT�~x���?��U���>�5�)�������jE��H�Hw������� ��VT`���A���{1��%#!��

�;�PyaBZ�y�#$l��ǥ����|>o���n�7��=�TU�(�3��y��Y��>�ȓD�.>�}3�T��a{5|���?�W�k,{��"54��M貗��|�nA��ۊD)հ�&H>���{*��2�y���d���X���ǃj��vHH���ԯ�REZ���6@����9�eM�`d�ߥ���J�܄�#��{��%m&oQ����������a$����Q;)���ne9 �����K�Z��RRw�k�n߲K �L�b ���w������<j�*���h�:`2���P{QR'lB$�C5?�W��r�-��7s�?H�V�I��^ �Zyrv�
�s���t�ԓ-:/q���P�o,��>��\�o%�� �+�u3j�|s��L��rX���]�-�"������Kl�X�-��r%R����W�̶��#�c-r
'p!��B�^G��Y�3�I���*��K�6���\��Ü�0��@y=E2���Z�W^�)a1-�t<b�f[��{$�Om�yѵ̭�*�J���mx'@A���f��2GSPmkR�L�$�C�P�Se��My �� 7%�|�P^]�����+ؔE@��Mb��ϣ-�G�m�vMW�5H�^0��\9���x>�&DG��B�&ƪ+)����M_��ĩ*�*A�{R'1�B�$��o0x�푇d�ѓL<�<���!�K�5#}Z����������
5��2�$�5'�3����5�KN�6Q~[�}�+��I�%{�����ヴfA��`��Y���zg)>�����h-Ԫ��;�ȗ�T�=7�w���#J \�i�ٌ��-�tԼt�j��Xe�frOE}#y�>+�*qa7�A-JV)���uX��,Ls�8��G:S���>�~W���~�y��U��ʗ>�7�ʨ�+���N0��_��GV=�}�處e�x��uFXl��<K��;�6�`��`s�W5Ѻy�r������������Ov�˦�Ebu�g 7��s2���h��(P�hT�%��f�׫4�����,�����|�8v�+}t���菔��V����	��7��}�@��
�����.�Dn`g��M����������ʭLp����8��"��QZä�̿���^�Ju����'ċ�$����S����Rj[����T����:��1�&�$�ʪvD���ɨ�.I(=!�=G�?`=SY'H��=a�zÀ�d$/˭Z�[xrRME4k([E�_�& �06<�5t �F���U�5L�^��ȟFRZcV]Z��,�h}w�,���)���2H�c �g�!���u
��|:�*�3�]��R��6�����6���>M�N�w鸗�`�C2�pawH;�r�Fc�nd�h�(�A[>U�OCS�!�@-����~�P `1%c�k�d�哚%��o&�i�lպ�O����Tb`�o_o2e#���a�5�8%]��5��l
��o���q�}�#���,�Qm`��S�jV�E>�jC�m��3���V�$� فvt���/0x���B{S\oz��(0�*v
��)��r7m�V;����m- (�rGg�Jƭ-]�O�q�%	�L�Hs�dH��μ�b�ԗ7[�c��̷;��zM����#�Wx1EV�*���6����x<��LS7k���5�C0��P��ٜ���=Bkr��k�+�_��qEu)�T�IW�-����X�wu���9
�����%���x@$���Ġn�w�5�1�i�08��S ����d������:� ^ts&� Pc���0��=S�)k����#S�P��*�b��j���R"�����R����>@�;��B��ͱ���}>��������)�]���D�.��R\��(����1�� �.��H|50t��B��[x�^ܑt?v�iu�)��z�kU�XX��%O�~y������ӓMD�C�_9�ʛ�@�V[b::
#���"�N`��Bh��3���mB��_�Y���-�J�#ϴ9#�Y9���2Ĺ�ɭڤ��V⍣5��B�t��':���D�Z$Vŕ��Ȳ]�e�U]�;��!k�yj�%+�Y�?���F��*ɥ�P�~l{(��;����٫�� 2�{m�[���M(��?�������@��K�ܐ���?�.����i *Iˋ%K�2�q�sK{Dթʇ�,0��,PG�3��c�o�!���[hE�@ŠvȆ��>��A^`�3���%l�-�͹x4���/��z���no���	Κ�5�y紱?q*��kJK����tpl��-���x�'C7�i!W�u�x�ܷ8uF@���䔮4���x��v'����M���=��&�ʝ�����#븼���x*���rG;�-P̔���a�
'�� x�O^��(��+�`���M
IpuC�k�C�ִl�&�倿�� �����@t��N
2�t;Nn������p,{-�T��ڵ�%�U��i��.�)n���]�q�����ϵ^P���`<��/?v&�EI�W#*K�>���g1Ȼ� ��v�n��Op$,f𲑏1Q����K�52֝��B�T¢jF��ϥ���19C��Q�#q8´,�y�� ;g�%M�␆��	V�="��4�-����7g�DA���Om�˕}�֮z����Ϩ\�$:�c �' ���c�GKK$��.VwJ�9�敲A��E�:Mm]�b �1Y���s�,p1M<�T�2T�F��Y'��W9G_Դ�b�
�w�����.J���<Q�T����z`�K�� ����,��N�����@l;5�s�Y��ڇf��e��*C�"��g��|�5,���ɣܝg��:m%q�1f�S[Kj���P�o��Mb ��DSE��V"M�F��J[|�d��.B�P�*.å������%K*-��2�?w�� aW���ڹ�h��� ������l��_6�JhF)grS�MQ�Ԗ���&�����2�c5��>M��Z/��x���B��� q��*�o��d]�O4K�[�=��{�o�i[��:-���g�!��W��gu�'�d�����(�9�,�� ���pU-����_�� �*=f���#���=����	�ܫ�pƧ~!!�;�]!�/`��EJ
3�
~�dS��dd6n�1���픝�&��HO��-�7M�&�
���~Y)2�¡��}�	#^o�`V3�<Fl��k�שޕ���A�vev�H���m-��`�-$�ұT�	�xp�!K�p *��,�\ A�ղ��'`d�K"�d	<��K����!�8D�B��ڙ|a_|�bϨg�y�l)��w$8����#Y=��^-����N�`N��'�L�F��~�#�4; -ŧ���k)L�
�h,p����U6Բ9a�V6�͞cr��5M%�k	n	�q���G��>�B��iB
�H�)�i�#���]�Q� ���/�@����"��}B�������sh��9���1Z�TU-�:�?��5C�劳哌���x�<.���JI��L��ۅ��"6�T��Pr�54��K��0�����a�H�aj�-E"O){C['O"�e����ɥ����N�t�
��Ǿ��޾���w7��i���z|Q����\���,��w�Q����fgV����,D	�A�������EkP� �_&�qmu��j����Z��h�Rk,m�T����m�����y��h�C��Y����?�x�M�-�p���Y��[U����G:W�:WU��k0���K�)��;�����7�����^JV��~@����$jw�I�+4�ur�3���mqU��0�SfL0T�}dFnmc��衿�H�u��<	��,�X�g��+�H�Rw�i�( �6G(F�qa�[�Ę`�{&y�%�o�3{�)�C[�*�~��2]c�K�H8@��Gl[m���A�O;���i�a͈����ӱ�opᾰcH�F�V�d�ɖ�����-�{���:�JX�^�d>�n���6�3�2d���>����+98c��5�~�=���V�Qyf-���̚Axt�m���>E_Vt=͚��t�t���0c�(�q]&2t&=EGL�jeRH�>Wq7\�f+uc B�Ffq�U���Wi/�?N�v ��\�o
۬�y�'=�߷n��g	m�{g�P-�8��)uq��8�E!~�d+'��,<��?��Y<1GY�U��h��`����yY͏c�W���G��x%�J���	N:�ue0����5��|�_�3�s�W��J�coyQ-�:y�=0�඘}W�i���]S�A�7LM��U�m�ᣗ��M_?��[`{.>},����ܒ�1�t��j]q��U�փ��v������C����NM:7�ggdG��~I�+��h�AX)�����BB-�~TXHgg�{����& ����)I����<$�ґN���B��@L�kԙO�C�"y-q&Y�u��h�x�vE}J�T�/�I���0�ů��ϝpz�v���&`���#O�ެ�0	ܣ��V
f~*�x��"�Rt;���d����W��K6��]_�^(�s��M�,o�5^�lFm�E��
ν6H�ʞ��>:�ڏ�+�l3�QC��e�v��B�}k���O��
�\]+��ӳ"�f�O�Ov��*�+�[�[S/=VxI-DDn��t�e�P�1��qe������ӱ���l�ݐ�Y?�mEn*J6������x�$�Vm�j�a�O�����n]�9j�R�VV@)�p~I�o8UC,D��:lƜz�-j�Q>��>]����
S�Wc�'��~�F��/�}�K�O7�ԣ^j��:��.�KAz�J)�KVp��pӚ#�%�����=GO���U�K�lN�c���*-� ��b�Oh�I^�&��ޣߑ�r��m�����6���P�T!f�BLj҅�*z!��`kj2���^c�_;r�x�P��RA�MQ)��k�i�����n���|�喸�aϑ��+�`�fYq=/)�R�hz��䚤�E4�_��I��(EA���KmD c���u�k�y���
]0�.����I1�J����n���&�,r��N�B�8i��Î}0��[�&�� �fL����� �Z��:ϼ�r��L��7�GY;e���������?WڰRc��.P�Zr�i��/�fC�`F	7#�/��F�i�_�z��0���#�	�R��M��F�̥`��r\j�2�x�t6R��8��b�6�rS&�?����?s1�4��ΆX���]ؑ:����G�ӂ��"AP�Kv���{x-��7��
�v�5��P��*�T��k����F�ۂ[=��E�aƭ9�hqފ�H)�`��&����
�3X��+�������zeփ���P�f�:7�H6>5)m�Z���"�"UL�5�����7���a{|H���[�/�ov�g䝷���:�\3�[u ��?T���n! *"�Kހ��Q��m ���� q�ע��d�����7��%j*?�X��﷚|�F?����.z�fN�k�$O���{���pvV`,	Q��	��Gt���e�*dd]��]ˡ�ÿWHSA=�1�h��eJ��,_��n��Z�E��$��G�&t�)��p���=��V����� �-��ŷ�2���}b�����81?���d�P��8tXP=pUy�����4/�@q;�/`��ȿ	�jC��@�I��Z�7�ç���lϱY�'e��Բx�ZN\��E!�-(1z���ծj�H�@������͘�r��z�W��9gf����Y69�69l��oz��f��H�^�m�-ך�G����
�}6�0>	w�z,��Gbʔ�C)ZGUZN,3S��|�^�;t\�*E����H���se��kY��3Ù�]w�}捔��>\Π��ӂ7r���:/q>5����=�^�_��l��74��=7�%�^�,��p���Mh���|��X�"���qd��[��&Z��ĒYa�K��(.����ճ�R������B�kŔx@ps�`��T�Ь$����uڋ���1�vJԱY��c� �J��=��v�~�ÂY�O����4ь�l���M�[�+��e?�M����'����S)*^���}�U�Y�^�l�2�aP�,�w%�w�\k
y�w)��I)s������$"��s
�[o<�A͡����1��,��O�\�9���Q�W3"�v�Ľq�S�����m+�����i��K�nV'q?���fF�_�i���i���T�ïe�T�C�u<3sL>�W{�%L��^HaZ�v�1n���(����t�Ѐ��g�u 	��*h���B�x�k���?�X�4#�L&>_� 7�%<�I� �Y=�ɥ�W��e���3�2�Ǆ��N$Y�&���b��Df%��1�UO�����j��f@6m�Rmt�x���O��::\�ئ|�D.¼�?V.�sq�����z.RAh���ȱ���}4a)�G-LU���ZL��m����"�"���Cb�J�I���E��9N��� ��:��BO�o�-��Q�98�ڧ�V�����Hg�/���_�a�����P���f{S� �r�fPG�������5���� ���vF��lpހӘ|d$ݛÃ)�E�Q�q˦ǲ��~̖j���4�s��������V���g_E�_��#����UUNW��t�)�ϱ���3�z���3^l�/���%s��;�N�����^#�MS:��0�����8r��*�汻 ����O�����n���䉫���T��1@�s�����|&�@��H	�6�%�Q��"w|���W��MirPw<Q��6"HF0�)����!�܊n���z��?(-����Ch�W�a��x�n���\���siO�v3�Q���pq���U
-Tb�![6�.�ŏ��L���Z�'	��qD�w�U�����i)�	�V��Tŏ��cE���mn�ĵ̞|�>*\t<t��u���K�w���IR��QOf�&M`k��mw�x�%�_"��Z���,���k��g6�����Q�T�EԽ�����XZ��s>�:�}���2&�����b�-G�o��$�E�>�@��Ӕ�li����Tda�l"#q�WM�='��9�v�I�
ת��s������E����7q����E/Xes@����%�VM��ڀ���e��k��Ǖ��,)Z��gL�G=|�\O#�입ZW(�.0��l�l��6*ʢ�U�����{�6����F&I�B�����,�0���+����9�G��?0�A��C�X1���m�h�{�:,"Ȥ��<�E�27{�O{�.{)=�wd09B\:�m�6Y#�p����	��M6 ԽȜ�7��V\78}�2�����y��>��tb��<*˱�a�T��Ee�5s�<'�����'��|3�h���y=N�3[f�e<�>8�5suլ�� ����F�9�-.�Q�7�𚯃 ����N���omu�N\g~�����Q���T? �/o�v)���q���c�N9���5�z��ꁮK�B�q]���ѩ��V��냃�EHM�0�z;��S��S�X�|w���Oߌ��a���s<����;!+
T@#ruo���2+'������,9��� �l��MM�m�6��u4.t��i���h`+��LP:|xKe���:a�ZQ&Q<�OÙp)gX��s,�R3�!g��S�*�X��r7��>������J�d(������ގ�[xB�S���C���@.`��V9]\�)��g1�B$H����vh�����l����a�)`K���}4sdE��f��0��"Q�Kx�����Nްz
�y�/����H��6T�L? @x�{'1=k#�3 h��|��� ʥuB�@+�Ԣ��CP��B�ˀ�Af�ho��!�yӳ_����C���J�J}o�t&xd��vi/:�1XO�&�?j�Vy�yo�'��d�s�����n�82>p
yG��\��Q�\HE���{��0������<�\�:&�U�\x�&,C��%ϣO������:�e��i��L>�ٮ�,,
�ÓŬ�Sv��D��8��`�?��x)�k57f?\^�|�1o-�1�^#*V�4c��y�&�d8��������3���̂�cO�������td�dwE�o�o�W�/��l������*)ARխ�r4#tC�NL�(!�:6���#k:(�3��}A� �)\|X�jь�F���T��;V�ϲ����{[Ut�ÐW�˒-�Ի�����g|2�İ���k�~<���Iy���a� F ��Z�s����i��|�	�0ޱo�)ܿ״4n����V�0�4��ǚA�/������rsu���a���P�?/����O�4[ˡ��;ͅ=?�=�Fwo�)77ē}%�0u��V�H�k�1��+�y�� Nց���`��	��'B!��.����s��vu
��;��w(�'>��������YIڍA�B��s��Uk�6�L���-ؙ2?AG��,R�R��'�J�7 ������D���D�M<��8��d������Ԅ�:?��Lܠ��t.� �0B���šntϞ��@��P�W�(�N��?�4Ħဘ5&�u��$Y>������ǀ���C�wN��x��4I�E�~v}7R�/f6d�c�.S׳5�4NH�Z6F�k�\.)���/�KӍ�䆄t����%�:�T�)�,��])%��{q����$1�T{����n��4���.<
�| �~ùNႯ6@�Q�.�n��X3.���-��\|Xf���-X��'HE�*[���~�n8=�ZM�X-����\x�$����2������'�BT`���t��.r-OJ�������I�>~?��Ϩ t�����1� ��,��cN3����������ҽ$>I�%S?�!��N�dA��*�Hr~��ф��T;fM6�3?�S�WnU���~	2�y��ʤ�/����j��J�4A���3���މ������c�4L��.���c�6��1��vO'�p��X�y�6&J/����4�hU�*��Q��t����1S�o3�=+cV?��q�qR��e��4joB���I
��`����o^Z�	���>6���q�J�BFQ*�A�{�œ�ٕm�]V����հmd��>Y�tG2���$#o0���0�UYPGp{��%�WE1V�t��?s;����1Q�N+ �2%c2l�ݝq�"���M�k�hJ����g��ZY��>�FU�P����>���#N���Ǧ�uJ�]uF��|��~�xd{��ܩ��/l��3Ա�9w�݋%�V{s\W�TO}�4̗�q��~�3�<���*j�Q��� ���.�rJ)���Y1���^�#�L�eȕ��t��A�϶4E�*���@�5�Um�<`�����>�<�� ��=�:�ɑӺ�TH��W�E0aP����v�������l�������07��|�L��$T��	D���n\0摍�ˢ����F��f�\�47�~<��>a������ּh.3�����6��j{C��-Q�q�a.���f�j���1;�*Q�]懁�ۻ}:)'�_Qs���c��������7-�:�Nm��@�ms��X�d9m�9���4
�Lu7]D�E#_����c8X�k��٪LC��ኳYèگ� ;Mm�K�$�;#���`����L�+*�A�<� �40�V3Kw�{e�����Lc�)U����0	��:;�;ZA�{�-�q�����t˸�G�*��f�X�D���d*~����K��g1Sx2������U3c���jV{�^��w�5v�`��gK��>"6��ze��RˈhW5�gGd�[_�Ya�V�`-�ru�=&�藨��^;��~�q���*j@v���g4�7����4�]��fr23j�5��@��`)��-��y�0'Vp\�6�xy�M	�[6F��1�y0�o�W��zTR28t���P\l[�9@��>+V��["�""��%E��P�f��ӊi�ڑ�ύ$��k��3�m`�]�V���ǧ�٤������洭oCF�9.C!7���T�Ɣ��[�l����2�7���\T�����(��^�.�w���N垗��lH��R�"XN�D�B!�����MN��6��&s���	�d�����3��
mX�sĩA�ݯ�n0��l�S�2��w��
55������X�3Jţ�r�"�Dh�X��k���{��%�&�q��̝��/�����5	ohV3b#�2�P�*���xe��Q��(k���I�� ��;D��-�̋��k�W}���k�]��J�EJ�T�8=��w�F#��W��9Z=B+�V/e@�A83��E��p&�
B�/p/�x�o}�!�H�#�K��q�G dە�)�H�w[�+o� ��4Ԋ� S�Ԋ���h�c�S�[�>��.%[�\=�M����dJ��ܖ��Ӟ�盤�[1E벡FO�H����uQf	���B�A�[�Gx�?FJk)��"}���-���i��*�'��9��)��F<���Ug"+�>���E?�o�TbMV�Ԉʰ?�k�!��Ahk�!�� p����`k%x�����D����vkiݚ�4_�emf�b�&�K�Ü~�|Si��;����9�5�ʄ�p��|.5"�q�L�a�g{�O���h��{soT,c}�O:��0�~����F�$[�ΟB��&T��d£�Fj�ec���'m�a2��%�p �!��Y�5H���S��hv��F���9��f,�5��j�֞���guAX�@�h��%�E�Iq�W���hAZ�h���iY(�v'}d$��_�g^w���e�9�j<�� ���[�鞭�f��Ur3r��s�M�h׵��8�%޺��8h]{����\�/&���]��`G˜��h ��D�U.����g営\"�8��$��a�/�S�M���W����p6�;�]LzV��l<��.�G[�P_�~����<-��A����.�'7A�_=!0�Iny&
)��J���7MA*���BZ�Ġ 6�d'�u������N=�k���T�7�W��)	��L���OF2A����e���$8Qp-�L��Y�i�XN{�̢/��A�%�+=����Ma�)Y�
Np���)��hՄ�Q*&�8�����|�G;$���Q7�Z��B���i��vRj���x��w�C�����ߥI�0�g��&�����;U����$V뽑�����]���U�+�[:|��!ڋ��5c��Ň��)���ps~J�arO}�\�3�tX;���~C��~yRL����K�/Űi�K�l�S/N��
���P��G��e6��h���pͣ�b�۟��A���t�2�azYc�{N�L(���L�w]��َ��]B�7.����G��c
oi�{$��+�;���c��~8�)�l�/j%�t:�B�h6�B<�uz{^f��\[
H5+	�� >-�4~��7�:~���N�@�pYkӤ����E.����,4D_�@�\fD��f�����ЃVBw=PZ� 
@5R�ہ�u��㖂,��i�B^#cDI}��#�c�, aUU?����ư\We��x���/����Ijl k&y:ڠ�N�)�g�[��plD*�sZH�ڷ�|c��"4�1�yg:|>��[|$���{��7�¾�K��	)��� O� 7Y*b$��� �R$p9(�sX����Z
�������'����k
�B�
ƭ�QjJsA�P��G2��|wWY侗�9�ݸ#�H��Z���w��o�C�"����ayj�݄�'��`���^�0Mcb��ӣN�aX�dE�R��?�i��**n��qm�����(Ec�:L��T����#��9	/2�ܧێOPI_>G��hAх*�Uw6ц�U:~�\ }�jd�xL�����K�c�2�,�$�p�Xʔ�5|���/K�u�9~{�c�5��@��9�8nr��b��V�+k�%#Bsr����A�p�
J���S����@�e�d�s؆[���U`Mr��.���րb���f��}��4qgpؙa�ޣ
x8yD��� ڰ���w�ہ���P����c�,OX�>�	�V�`v����&�fo�cO�	���'
.Lw[sM^7�s������#	h&"^��^
W
1c�Isp��[�v�9��ε����-i{CF�v��Lb3��sc/�;<SJ��T�-���?�����?�����|����N�:?k�QΏ��UAE�K�~�b_C�`X�l�$�ڦ���q4���"Ld�P��3�#����x�RO���y����C�҃�i��W�{o�SDM,w�����8�?�}y�9~c���)rNp�QK3����>W�rU.��º
.�O�h,��f��91�W��wK�vt~N���H�#ª��q����}�:9�ƪ���x�	��Y꽋6�t�w��h�|�̉sF�r�$��
���9�JUxh�7�"�?j��03�F�!vO##2�>�b�"s�0)�����00b�5�ߘ�e�t�	���4$�N6��L�~A��_lՀ��ȎU�KG�P?�,hd��Փ��b�޸_!2�Mp�h���H���+�v��b�.�8E��)7_��`�O!��@@�՚%D9a9a���A�� }�}�M3I�n�'��}N��ɔ�&+P9�c�R����˯�����@��&��铷R�;�t���Hm�?�V-w�����UL�'K?��Q���S=�-n�ǵ����S���tx��3/TLEm�j6�gk����x��P�C~�Ŋ��E�]:���&�7��p)9%H�=�����LvN ����y����H5�+3����F	{�6���H�hʂ��>~��ўDl�B1c�g�C�ј;( �V�[ 7�Ջ���ϭ��%���6g��f�������|�(����&%pFN'�ʕ��K�T-�����3�pe9��J�i`JJ�0!�$S۲�ǁ�8���*�W:b�v���ju��ߟ#�9��ۂ064��T ��<����s�4�a�N����F&��ƾUO�Uļ*�ރ�: c-~�ɠ���%U�9NiߩaY�ï�&�ޒ*�z`�h�P��"&�s �ݐN,PV�M�}28��b����A� �!�9��I�Q�E,n��"�����3<wIX�\CغB ��X��7���-�H��L��G�r�닳���;,ME�!>}���=�[��,��P��챺,�Aw�M�%��GgU{[ػ�o�8���K:�ޏ-D��mU��>C'��vm{��R���$�w%!7��H�?M�1�,������G2we�o����M��ye��0������u�)��An�1l�^I��G82��ߖ��l������Wv=�H_o��!67{{0~t><��Χ;/�bn�6�R��S�O���NMV�V&�-�Ă-DZ|��K�Jϔ�[��3�n����6��b�Jհ��R)�;����E. ?d�Ӂ����	�㖡1v���V�b³�v���9�S4uJ�M��S-ND���1f�_�X������k����+����o9��WZ�c�G);��.U�C:�yވ=!��b���.M���,�ځL�f�_���׬�z��f�n	���Bsf���aorb��`Oi��? ��I��[�!V��&��fWt���#�R?��򥔔�*]r����DM:��~�����t����f4���.�ɭʗiq�]Ƕl���F�/���_3��+�߅ ��r!�a���N���6.��'g��-�	4�j8�޾dX�ܝP�hʶ���o+J��*_�k"���r�Y�F�>�1���S��wZ��O�H��>�(eUSB�̕�o�y3Ǔe�f8�v^ 2���g@N@ܒ��.�\��kDC,ZË�Eͷi��c;���ĥ(�|��h�����	��6 ����2���j�r�ߡ����
� ]�o����p�Z�Ε�Sv�{�������G�k���jry4����T��W�.���P���f�%�L���:D-̳�b��w��Mg77y:�aǭ�c{c�|�3�I�!p1�sWK#��f�"���To�������<��zI�����t�)���#�iP2�Ӯ�VVĳ�ц��:t[]H�R�S�J�i
��@�j�wLd�ʹ�x�(��I�c�@io�O}��������~1��z�=�qى�� ������:�*S<���W|R�R�=dm��9�/�x�,��S�L�����F[? ��d^��p�xt�Ԥ���4�wC.���&M��0������Ϗ�SL0{���4�����7�M�-}p�NZ"�0%
��+^(��c��c��O.�<�vm�!������e}[�>�S?:��oX�㋶7�t#l�t8�gä �7��6��D���N�B��rs�h:��n�ZXM�NR�?�g'��.�φM����p����ج��m�ꋣ��dt�gc����(��o�l�v1����w�e��:x��+x\�Dg��^m-[8R�'��uVW�G�q�.�E�Uw��<�C��z9�������5��`�Y-��j���B)5T�	�WX{�4dQ[�:ĥa��q�?VZ
]}Eե-�P;ΞX�,~����ȶ��)�!�:�D/���ԓ��H���T���0������|�'VuQt�m]�ܐ �qaʘ���~�^c��v����[�PMgV��h�Α�zR{]t]�i-8M��%9�B6@4�(�*9��O\��~��L��.	�"0*�V�6S~\�j-kH��>E�N�����D�-�܈�!Xg1�ƞߎUV�E[�#��?l�ZIrZ��4�&���M^��t�Sʇ_[`T��V������JO��ɒ�苻a����A��y~�l~6�i�M�P3��/#��uC�ّ�2��[r@�З+��l��:`�F���Y��a>���Y�J?�x��2�/���8���G�ȉ~���P� {��q�����\�����,v!�����	'B2p�S
���#D�y� �+3n��e�yC�V`���Ϧmlro��}�Zrd!����m�G�ly+��Ԏ��Q��<����'��1�Z_��<P�@H���0�f�a �ƴ���<��umm�8��9w.������2Rm��|�KGIO���Q����,ǉiM��]$僧`�Oo�������T�@��)�$�(>6���s���Cj���ylBS�u�;ՠ�
{v��_�����ߤ��!` ��!B��wq��))$G�@�C)��)Y�ii!R+%��fnMت��e�|�0���ح�����ue+���>�6 0�:e��o.R�20~Ug.�NP�S�l�R�It>&�(mAJ)E�Z�`��>�73�:��z���<���pN7�m Nc��w
?r�8�<����h-Y[�Já;{ە�be�+� �7/�]_�·d/��c��6�0�9C�n�#��m�"�K(�lpx]�l�MB���>q#��#���VE�G��6{ą���`V��@N:zW�e����8�.ul0=���s���7��aP~7�����rv��*f�d)�-r���ל��Z6~�Zn�����R��]��~�����y�jx�\}��Y��a(S?u��zc֔5S���k����C�lXR�]}����FIr⣀r"�:�f�H����l�A)�Y�l,���0�nQ����s��845�F�� �em�OgP���uC�6�V;�<`�aHr�*wR˹zD���b�3�=����}x�� @������N�M�j��Xտ�VC?�I�ZY�a�b�z]�8%�2ܦ�7^4a�p�z�H��0��/�����ǚkj0�/���t~���1i6�)Cu�!���1�'h�P*4��ZH�n|�_�"gq�n#�1��aS@oq�R���IEB d	�+'I��� ��|�'�������X�	9Gx�6ˮ��D���_� Nd�"z��������~��4�3����6{"c$L��y����>.����9��G�$����8���k�2�v�~���4R�Z�5�p��~K��[m��V���kS6�`��9f���m#���K��ڞu���T��hX&<�$���^��Ҵ��~ܽ�opf �y'�5�y�G�dm4��@�ӄV��_"�B�o�3��5�,ǫ�sL'�1�l�g�+A��bW�~����jh��M:5
�a���3?�5�7�TM��������#o���
�����b�Qw�}����T�փ6g�g�Pǥ�N*�5�P��`	�`a<��Lx��l4{�H7ùN(˿�zr�X@] ��fP�f����*ܢ����RW�����#W��u9L%r2$��ԛ��=����=��󟕨_t���� v�P�ڄC�����Z�����{/���1%M����Iѱx%S��:欞��G) ��������{�����xK���|����8��@�~�}�L5�Q��]v�9�@.T8�0%�{Q�Q�NE
>���(��3N���;��8[O����j�y��.=c��+�oAIԽɷB�@�'�a3�D:�7�T��d�B�u?I?T��n��ϒl�}Y
��*/�ji�t��U�Y ����@�,[,%t8�=1s��+Dx�i;۶�\���=�p�\.&�yr\�E%Y*OJ#��˃���׵
��w;k��1�	�,���3b�[�)��j��k�2%�����0��2.����'l<���4�S��R�
Q���荂"����U��^��0�����`�uT�ܤ͑M6����9c1�ɺY>0���O%eW?�'�2V-�زQz�����������}����5��>��Y�f�4���b���52��9%��(о�߮�L���U)%F��$�	���:݃���?�y�N��ӧY����;"��\J��]�pV�O��$���(lF�,�Ŀ� ��Lc'z�x�����Cz���ox�8�w,���~������|X��HC�怌�y]T5{�Lf���6x�4/�N�/�N7���U��ɋO�1�a�l.��L�-����'s�Q���ݳ��&J_�$ A?c�FB�$��� ��l��S��&<�8qh��b�$l@�w���-�g�̯���t�	��=)3-=�p蕺�ǔls�����E��/i��
V��%5e4��8~���x�:\�Σ������lL�� zg�\g$��n[<�֊}v�*'��J2f���cd	��R ���Sk��BN�[kǶ~�L�Y�(ϭ�����}�dÕ|���4鄃g`3����.v�}��F�k�N�y'�T��d�&��5��w5�m�o����C�{'���m;]��>���'+���2,8,�&<�&$��߱�!��%d�����I�VC�(p����A �d��ڄvT0��Kq�=ϕm���6�;��	�_�=�n�\03��v�x�6����k�1-4�BV�`]��wU.���Q�e�C���*f㴴�U=��s����[#^z�;�j4������IK�������2�\FQ�#�Ə9��Ϛ�R䏃�`4�;Bm�3'�������W���A:Yk�s� �{�%�~��:����{�p v[1�WS4f�`�<-,ۢ�#���vV�*sІ�MʡZ��R��Fn�9g�O&�z�zS� }DS�YY(�����id�B��<�m|;_!�N�_���=���I����H�&�p$q^S�P��.B�K$Eϖ���zr�?Yy��~�_�*x�������S�b�_��(���*[�P@6N����^���,$@��yA�����q̽
�08LN�6a��i"r��6Òhc&	�쇂R��/#}�UF�Y�t/"���W���|�d-o�^I=�8f⴦9ۙe���7j9��~��Wv���z���P�S��[��'�0�o��5�#�@zИ�W]Q��JJH�%�p�-���V.O��&N�v؀��V+^KvJ�%`	�a��V��ws:Ч�AsM(�;7Cٽ��������S6�Ֆ�q�3c۴@���#K?�(k"�G|����$��G�����zIU@��"GpWn���~Iƥ�T�'�H&��񹢋��_�W_׷LA:Ce�d\�k���D�����<���t�W��A֝��� s��x�=���tjی��ʓT^�y�e�W>���fX�o�b+~�A�ʥ�ë��ى��@�d�~�z`S�!������:刣(����3"|���Y.9����:f>^������=gd�ޟ�/�ʯ&�I����D�3�q&�6V��	36Q��";��Z����K3Zջ��w��b/��ݩ��R_4�J���e]�h�Q�A�$���µ�[�:�B)!�v]�qkf���
�GCE����:�ћ�� VS䓴|��p]��[��];�0HW����0��i�n��������w��g�Î���2w���Q��m}ctu�f��#Ie�{�4�M����|\�&�k� ��z4��tKO�^�i@[�wJU�G׀�mx*�dr"RMu��?`Q#�q�aS������Y$�жu�n�e���>��wX�ˉf�<��Dyt9�ފ�#U�s ͷ�m��y�Ѽ��,�ލ��IR��o�A��QX�C��O���m��}��jT:���ng�͉�:���d늷BK*�c�;<���Se�q%Hn>#�����Z�nQ4�ʔZb�8����&u���*Dk�#N��Qu��r/�o.�,R�l�&�k�����}�� ��=�
t6�|��,g�Dp(�	���D�@�y�� ��"���!C �r��n�C�{��:�����y
�:V����闳��鱾#������	�A�E�(��� �VY���]����#�ϝ��@�� ��L[p�vw��]rd�l�ےd��>��b��@yZ�pr��ژut
%0�g�]E����^��do2(���ȅ_�n�E�hh�[,����� 猚�e�~,�(�5:,�ߕ��Lx�uH�q�	��%.~6;B�,���������&[�5�Ġɥ��oJ��F��'�b�����!L�_�1���D0Vl�8�"�A���)K�o���ϑ��� ��+��N'/���̄M�৉|i���.͵��n߅�?^�{�[=�M�� ��Ҡ�w�r���;R�V�. JP%��	�Jż�V�ԂB�]Y8�C������8�%yg{E��	�mx� m�b%L�G���w�ʹ����e���eor�%9�,:��m�E-��On|���1�W��)򜳱�e!����U�>��y}�w�H�i:+����S`���L>���}�eu��7W|�9����8�6gA���������a,sy�Cx���	l���/��U��{P�!P}W�E]���$��u�@TH��^v�͛�DB��R�|{!W������j���s�|�@}>��(����'���)���S7�7��$(	�w3#�x�R��;y�S�廵��7�%d(+�a^CX6'�4��=��XеKr�G+	%�F۫����i�O�Z��_J��%EF);i9��e����{u�c�E8r6٬@DSV=���M���#R����|@3��Q��{����~��p_���(�l&Ʋa��5�5�b7��F� ��L�x[�^<7<���81�M�K,�x�Ƅw�� ��Y���*�&�ʹ~�U�Q�%F���*�k��+��\6��)ݼЛ�LIf�[���!ʆW*+o��@RDAzwP�h�xb���ɲ�6�ihu�����iVh���!���?Z���2�y�6(w�������F����DnLNO��B/ڲR�����-� ��6�-��4BAI��[_?�B̔Q!I�*AKhM�e�5L��P�ް�b�n���wYۖ�:�9�{����ؾҌ�bSo�DNzY�_�ݖ�CT�}��ڲZ��*Dj�n��VO�ҼTꍯ�EA�Sܬ���[��I9��l';�j5�]���ww]���c1�����Ղ���	O%����Ȥ�|�Ʉ��z���c�������4�JJ��8A�¨��=H{�iDwJ"�����G�:��3@����tR����{�u�g)硸w&Q<5(Jq��}_T�n9�~���V��#)�Fu�ph�c�a�譯��Rb/Q�$ �ٖ H�fhE�a*+r�L$R�Q45�tqޏ���t�U�ɵ���+[��b����k��7��״XO�6x)���KYМ�x�9t绀�p��^,~�D��z��"�#!�Q=�{��`�j��n����G��~��L�j�a�L��d���/�p�QK3֋�E�|���!��
 ]������	1���ry��W"�<>�/-_d>j�|�ͯձ��c��;�.zG�����j~����ۣ�����Z�-�m�&��%_Q4J������80���5O�=F.@3�qWEO���������5��m2�M���1�2^6Y0_��;���Q�H=�G9������Ycsf-�C;[� ��-t�ۑv��Rd/��y-:�
9����w^=D�7"J�N\50�t��UY�(R�A�Fm�����=�L�?�s��R�B#r}����������\< &�.�Oǿ���	M B�=J�z���\]ܺ{qR���{6؜&�9A'��uѷ�@ÞO�47��O�΍�����Afi��A�㐚�r�.|4dw��+�R���X}3����� 6\P��{�U���6��7^��x�¶
e��v�#%b������@����ʄ�(��>[�}D,�>/�F�%��$~e�Bf��Q�(Y�4Gí�����0�m�%�����P2��>�U�v�Q=ަ�wX�bJs���S=�y�4n�����a޼?Ya��S�P3u�}�\QY����$7�`W9�4DA�	�Q�6�K�]�A���MFQM�) �u(�A�Y�&h&js3]��jPpk���2y�LJ��gL�\k�]P��DH�I�a]��'c��<@����n���Ւ>4j�rԚ��FR�<�s���y�c�\(��	�C�KR�H�)��<h�9'%Đd�2�ו�Xٖɣ���n�k���).��C}�LB:������rf����l(�p�;�?�8���祔�Fê�?L�aDY�x�����4#IS��jn� ԻNMlzFaI�b��C�����1��x������ؗU���O�'ܻo@�}ɟ�k� �����2�f,� �ﯫE�&��w:�X�������4�j/(9�W�!)^h=2�p9�����iR��mwo_�Z2� ;\,��?;��#x#�����ꁏ�$SikPX*u*����7EO��FU�X��=�/�C�O�);�B�6H��bC�=�`�M�e�f���	j3�D���P��!���x.���k^7�W`�Yh�N��2�Y��$T��?��FN�_����K��WT���a�O��w��H�hC�r����[�����ﮰ���� U$��g����AB�2D�5����4�Y�t�J�cW��������X�J�'���8������qyz{�H�N�����u��U�S�lb�!i�;j#`��2
^�;�>�Ї��DZ�@��22J��)+k[�OF��gA�Z6�HT��|�d"����LT���7Q�*��sj-8y�A�/���t����#�/��I��4�W�X"�REU��b=QF~������*\��G�3}��[�>�6Ò���wm��J�X�G�C���S�qV>�>��R���O�3a��֢<N�L"*���t�[���%m��ܽ��3���F���vDc�fl�@ʣ�0b�3xN�[��~�N5H��L�A�KZ�ɰb�~Vt�<��LY6q�J�p�C���9�Pf���ԭ�.���X���$m�^�X�ʺ�y�8]���nx\|�+j�'�t^�aq-�eeYsXپ���������H�݊�މi�� E�p�����^I��G�)^!LUB�ɲQ�E� �8-��j�P!���Q9P���^�w�*��u�]#���+{�;�2�`[�h��C;��_�&�����`#����T�����R�A����-Y/MPE~*.d������9��
٩G�����J��\؍�MЅ琔�	E
��`�*��FB|k�ᖏ��Lk�K8L��!�g�n��/��N �I��_M��z��3�-��!-%Pd�ՁH�����O���|cON���k��ܣ�B=@?ڀ��C�@TF�t'�}����a�C;��^�2���E�u���W]ݎn�$�D0����ܻ֨����v������y�G��X����j豈r�h\|��X���~׽��ICW]��J-�w+�#U�	<����l�!� �hx�Lk��Z]�ȜEl�f���!`�!�*�#��AW���A��"LY�R��i=o4m�ޓ��	qS,$:��l��K��0�%��F�z�䞏1'MbG �j��-q_�t����w,+�\Γ�0�G��6���$J�x�1b�+^��T��DF|S����&���?#��{,4uwU���z�.*�'0z�������aaN���<�_�"��������N������R���:����$�pX���g��m���7mߓ��+���*�\x�\����p�d�@iϋ2ou���ښD%1��^3z4��g2�GVݣ�/.�������.
9��L�����rU�A�{6E�e���r��i�r� ��)��ʶ��U:�n�U/��L�F�%����ʃw�;�����c�8��n�ן�C%�˩*��l� �;� @Q�q@"E����T܃�Zy�qE�1i��8�<��*�c��|��zdI3�iem���,\��Ph*��{�=��p7۟cD�҈	/���ؑZ�@rq��l������\MF�HۨЬ٬{���i�����59�^I�G:�Jߔ]t�w��u�:�c����;K: Rx�t�(��=�ސ����i$�~S��&�\�T��� ��V��0.7��� F���]|ߠiDA�\op�l��U��꘼��M���?1a�l����U]�m�gN�š;)�Y�-L�To�cn�P�����Kq��$��r�5�!�j�?+��o��6�Me)P;FN����hR���R�);�{FҘА�+��Ɣ��k�S����c��s��:~?�!�ؽ)��l�4&t�̅�� 	�E��|�agʠ���
�������2��jE�a��Hs���5e��B��2�V�+"7_�4,��߿#|�,lO��<=W�gMP���V���ׂz��6�RU��$3��E�|��X��b"�WN���;u	;
�û=�w[X�2�`��hg(�Rj�%���̰���$���y�a�����+�/��<�=���,N{WA�{�s��ϤP>Z�����9���3���Q�wP�F'�����A^$�=0�f�/hv������8���B���o��H����B����b2�+���-kf���z�X:�ig��L���g�������k(��S�3����]���XJT,o�?4����(�o�r���:�z-�
q��Y�K��DW��E;��px�#�V�^���fxl�[3V�����,��'��稭Wj(|e\8�7�3��>�M�*|�^s7��l[��"�	]�g����`�v
п7�zr3�1O܇ߌ�ڎ�t��7�!lF&�p��"1�����Ф�o��� �#����a���Io�$���/`į0����a���%a���̠~�#,�/��>��^;FÈs��凧�bB\�Eg�c����Sp~���wyț%�3uY��e��i;AUi������M���<��x����kkr�kh�o��g��\�R�R�P�䓾P��HO�z+p-��%�؝���A#X^�׼H�q,՞�&��T�
uc�Va��ܪ�[��#x[Mĝ�:�P�P�?!)V���_��MW>$��Vc~S5[Q�������9n{�j�$W #W�ğ؏�;�x8_:J<�s���|�7����@�A2Md���c^��T�1M6x�H&r�4�2O�!�?n�&;|�:,6-X+Qe"���͢��'���1��'��2�풶.��b�bj<o�~��t.�b͎v�F�nc�+�����9� ��F&�/I��>[�4/���$؅ov�������N]F&:��3�1!��2��1.���f�?o��
�~o��l�_xv\��e�w�|;�)��S�+I��C��-G"�R��u֌�s��Y͂=��K��!=n)����<���^�wP��R�k��z�ZΏ0.�+�3Ǌϓ�����]�\?�sv3w����E>���Q/A��5��O�� *tM��Ԙ�z-)��zH15V���0�Q&����k��ml ٻ'o�k�s����Oh&t����ىG1�u�+4&�h�/�o��Q[x�1�V�r5�C�T�T�i���,D̬�=�g�}oX[���%G�]�`�y9cP)�)N�@���� �gؑb}�3FC�(���vV
�*��e9�[�u���}��9�pL0p9�?h@;q�#�P��ٚ9qڙ6���K�"hc�ziH�9����������"��<,���e�D���fr�� (1��M ��B!����j�U��Bxp؅�!�k��`��_,�� �~���䒲m�H\��\Caa�U:8+1�w�\Yq^$��߾諉� 4����"\�&[�Y~jL��6��
���?C�Ix>?�K��>�&���!C}[�����U�{�w���x�.�#���g�T�/�Ȳ2l�؟ߏ���>W=�����4�P��٫��8����̴���c�
X�B��&]9�eF��Vt]5,��]��D��#n{iU9d5�R����e��	5�f��W�
���?C݋7d,�wSjsu��H�{�Z)�gW*<�3���߉7_&��`Soe3�>���+�~�+TW���R�AW$R%���ȋ3����`|�1�j��7L�����W�}�Ј���I�1p�Y�K����o��¡[����Nyv�J�>r��P?i;c��P̀%�Р5y=����Ĥ/?�,ݰH��c74h�A}���z
�c���F�=�6W�v�3x��O�V��DǓ&���pOЪ��a
�b�1�u't��1��ޒ��%(���CW���@��
�Z~�!R%I�~�H��-v5E��]v�m��ƤpN��}��""N�B6�a1@��px���gC(v�/T�	&��^%m��,�[��|�J�g0z�R��k�&�j��l��d]ߵ
&�xr���R��`����1��$����ǣ!q�io��=�`��g�5�;�Lo�L�9�Zb�]L��5Dj�G����أ"jy �2y���ϰ�����*���W�Q�SN�T�ͷZ��3]�	1�j����}�-O�����j5i�b��!��M1��W�10n�&�������	�?�����~����a�@μ����s�K�]��cNߵ��9�h�@�ɪ�n�?S%H����}T�����%����c�ooc+cֿT�K�"�4I���+ㆢ�l�����`-���]��6��D/���~^�d�B<ql�)�&����*6~�^[["u4$���`�_�$�y�\\���vl=нS����`m�����) ��� ����}�)�|+����2��p��f��L��б�5Ly���e2��:�;�o0�ñ���e�|*�x�t2K]�?*c>;ǳ�u3�c.Y+�n63T=>�T��'�Nr	n�UhZ�sU��	L���+gMG1FT8��9�M�&n�Y�Vu.Rg���W8n����:����
���+��Щd�>#�
)�n�X7�*O�`��G�X�Z��~Z��3�PѶ�4�N3�MR��=
 �� ���/�]ew$̀ �p5Y�O���Y���?��y~k�cL(���G�IZ�k�/7���2r�����s�.�~�n���J�𠈂� ��f
	��-��쬫h�3��G}�u�=,sY.���w�*��r�`�L�'͠-ܹFo8�	�D���dr���y���Jy����]��N�� M2��fXA��I�5%6�U-�D�;�_���PT��F4(���NZ���#sD�p��jX�=P�'���.z����q�G0<�����	pk�4ܲ,'����G�d���9����3���}Ix�C�U�Zw�;疳�/�v=��<�4'����n�)�0g	8Z��u�_��_����LN]ݟt�@�����ïF�e�UV#U��v~xF��5��*'�?y""�oc�O�k [�����m2����`R�jHP8�������Dl�xz�[Jj?)
�+1�3BI?�U���Y��4�(�^>/��RA;��c��$c"&O��	Ffl�����ڥ���>��߭�q	P��3�g��! �@S��V#�Y�Ѣ�)�0���<�!��rK�,�����i*�*W}�K-�D��L���8�0�[C�P�M�#'�6��+$�((��Ch�6J!�����z����-��)j��>�SaU�BڑT�yK;��q;3��D"���0�
�ۈ�}�v[�S�hE�{@�3�-$T�S��ή�r
4�E�8afv��ЃU�9/��{M�Z8�V��D��-ح��|�'�M�IQ*�0�"n��!E���چ��3�����2�d��En�-���1
p\N"�����=�3�X۝�@�bh�t���|	�o�"9$����H8�h�*V�����v"����;O�&�E��Dd?���$�Ă���`�N��0�3��?�
f��~i�y��U���4B�X�3����+`6>�{��{V���/j?/c} �|��M�y��T8#z�aa/��B��紉UK�G�oQ�)r�!��� �W�}�L��>y:k1����:;��.Fo��q�޹�<��t�  �fi
�<��&d՘�kR|����e_�O��`䩮|���Kr�g�bS{lX�n����S�X�o��&jV�bt�۴�ڶh=��ST��L!�L��� _���v�t�3�Jꕃ�'cG���Lo�f�g�F2�N�/'-溯�^�	%�'n��V��+hB6�?�k��zk�B����Y������\���D���^����*���ã�\��jV�!��썹���anOʸW�8���;G'(J�����"gN�;�>Z�~
9&��9h.��P�Mk����H#XF�\(�ӑ�lI�\/��SR�l]Y��`�|H��,|��T#�υ)ޏ��o���|UF|_Jc��vG�G0?|͐t�}LU�D�i�	l�#�y�&�jBL�W��-�?����*+��*��ͽ�����B����u�?kD=�H�ʄ�@�%�0ĭk��RJB`��$���s��x/w��AТB�r3}�5�S�4������a/���U"�"lk��D���tI>
{���ad?���< �C����z�{��2J�sÞc2'�vTjJ������U=�w,��e�\`���A����W14���=�C-����sK�*�֕˶5�ux��)�7����YVc��v��bc��,Z͇�R�츛q/E!I'U� �ߝ���u�C�m�w�X:��ߍH���;B��Bz�BS���.k�HlB?��"2���5�YpۘE)���* �� �<��<�GqԚ1F$W_G��=j���6�5D��(^��m%ć��ֻ,m�|pCx�����l{а�a�[���V�i%���4=߮1ǯ"�̼l�3M����B���';�uM����(��q&����bB���\�L0��x"(؈���^��G)�|p#~wH�.���s��^pz�x��HE�:���;��H���%�I�a��_]��Qm�1^{u?r�G��Kq�Qv�C��+�f�6w'<���1a��:��{g��wSV�6�e)����#e��n�X���C�H�'�>Y1u�fK�0���	J��)���ģ�v=1����0+�;��� �-��|�4��	,)� �C�1�[���S�42S�wX53�.�*G4��c.�5v�KAΌªo����y��X�/��X�$q��U�T_����x������~�`�+�dh�89��GP4����9 ;>ڠ�B��}\���,��f��I�_Xצs�}�#YWe�% �w�K�{�]��K򇁹���\�
V����3�z.%�S���&����cP���h��7����i�E������e����C��l�b����J��3�Y�|_Y����x�y��jO���\0 �Bnr59���g�����������n�&�?�͗9mΣ"ߵ�n�!J�|�f�H⛈����!,� C�����������>�i�x`����������t.|柕#�>����D�U%�����$��W��#�EPW�Gq���xbQM��hs"��`۠df��O���w�u'm�]n��t|;��GR4��.�벶���	qӚi��60��3I<��R��@�����*���#)رяe�^�ߓ��n�0dzʪ��--h�U�7PG��u�}:��B.�n��U��{R)��?�Q+<�;�Ԛ1�3��䦈�� �A���W~���}�^F����+tq�EPS�x��XO���P
8P��j�.�����J�����ҧ��#<D��%�[T����|���ȭ� ?��F3
+)�L��C���J0N4��M����GtE�9�o6[���l>C>���!wQ{3���:��^JZj���Ĉ~J��S�$5z������1��ǎT�s�=u�l7؞�=#T��o5��6g��9�x��.��K�m�P�hc)�#���5�tgp��'X҂���xj�
�<�������ΤU`rKZ�@n��f�;����\[�y��L�j���^��=dď� ��v������6yVl����Sʓ:�~4��c�T%��
zV��G8��E�~�,�^�p08z��cYxŷ����~��$3TP�4��{{��^?�OOa�eM��.��C��1�T[��
��A�K,�P����:|�9�����,�LD�� ����eSޑy�������DFۑA��O�0K�sO'�6�s������9mdt:D��0�Zle>��*�!��"�ʦ4�.G���=�&�,�q�wD�X��Ϻ���RK��Z���;��3��悂�$*C�fV�G�!�ޮqPT��7��Y{�
������ޢx�fx�a��?b�%?��$�
$�y�xA�]^a�Z�����_��i�U��P��|YX����G-�((�b۱t�K|���#�8̤fP�/Y���6����-W�sq��+_6�{�����W��M0�(�ķ�����\�ׯ#�Y�a=HW�pKT��tS��j&9�7l�H�z6s�4�&x�QM3��~IF۩y�����Ǡ�$å#Q�ν��Z�B��A�p����/�>��s��l}�+���x�|�H���+�8(�8`�Zq$���]�%z��o,p��2��)_::w"��aDi��!�S��o=��g��� ��)�A`��P�O���A� (_��n��<�5:�C�.�4�a9(!��5��i��ѥ���y]�MSV.���,`�]<��b��@`,����M	�d�$S������;�O���)��ǌr0A��
;^diAs^�0�<u����b�S|^[a���:��z��պ�:c<�{��̩C����[�c�����3ê)���v�TH�#�;��<��:U�H�8���`���ήc�M��u1�Y��@�B�j?k��S���1F_J�q�ڪI��hrƿ�/���}�޴��o��������uC7�����	4ɓ���7�������Y��j	Y'
�.ح��0��T��ӍT���4�$�{�sqDq(������X ����iJM:���J���[���-��X�ק����ΜA�̃xf�J���X�#�㊆� �.���P�Z%{.�7PW�N���(bǣ�D�'���>
j�W�10K�X*��$���v�<|�N����yY%���x���{��W�!hH�p�J�de���a��R��.Q�$F���.��B	��� ���+�m�ct�e�^�N���j���CR��֚0�~$�Q9�Ə�H��O�'B���5��M"�R� ��+��KE��j�j�Xi[����l�9͋�B����X�R�>b�m��b�Y@���mC0w����y��ᓂV�p�IA�����h��<��d0oY0�!y��Q�VP�h	���m�<�����m(w6y�:����'�o���N��3�tnp���έMNP�\=Z#K�m��ɛ�t�ި���&�Q��ZK0���W��c8H�S�(�(��� �*��<n�x���?�v��>�v�V$�����p�>����z����&%�8�U_XL�gt�`�Ԯ3��
���*𘰁pz�I�g�w��ل)e���f�6��e���[=���,��g����g;%rX<ɟ��RLI�(7���1rh�Ӵ�� ����w��0��D�5C�����i}�.n>����{ x�J	G�Osx.�h���=���!#�Q�,��I�b����π��E4�|�E(N{2iYГfp)IkE��e*}=�^���͘Q� 'P�<��(�����cgh��~O=O�2�qE��]���h*0�+�h=a�e�6	�~�dWSM��qo ���� �ca�j^�7[_���d��(����&�;W��j�f���K�C�^(C1߽�:��a�Y�mD��q�0��`BIw;�_�X����R]��1
Β��j���T���J�m�e��cC��\��MK�K�}n��PVnF$�07�;ox���T�j|{��̸�%v�Rݢ�*4/Q��_dpɓ�<�$�����a�a4~0�-�	�	q�|�$�K3	9qy�"jF����!��M�M��7�s��P��^B�#m��lPX��u�#@}��=MK%k*��A��t��o1����q[�ma]�I�{$ts1<�ϐ�U�*�1_�&ΊF�fL�G�c�ث@F+s$d��Mq-$qoۧ��61�!� �B
��r���`�󥼭���.C�b@L�(��+����@�P��N+͗�m��69�*
!����u��-������������n*~�8K��nPΘ��б|6�������9����9^Y2�y��ߙΝ��w�R2҅�@sW
���PF���*mwͪ)��z� ��x���MĢ'�������g��3� T�
L7U�~v�WM�b��g*cey�sMⅣW����\,@[�����8���E>���u������ �8V��9r��ߣ�p1�n�\�ˌ8)OϑT򑴿Cycy�~
Ř<D�q,"�<PL�Btź�7�pkF���@a�Ϊ�_t~���0Q���SZ�I!����@AƆ���� bI]T��-��l��5����m{U�z����N�.}��G�ކHt�3�%!�?�܎_���2̄]��-�Yt��-k��%L̗ӱ���?ao�O$?��Q$7�XLB�!Z��Ўim23�3])�TT�fk����#�B���a��-����(7��Q0����� ���%p�/u�i���
�8t]k��#F&p��6���aL�����m�!�[P�,uo�]S�P�%�˼��̎.Z]-8����G��&5BR�dv<Og�X��㚀.��3��]����u���v��M�6y�np����A=���iX<�nL�@s�2y]=��|}�yL�|�$�������
�,M/E�{zzP����}��9DA��Hpo'��w�7���N�̧�V�\.�T�c���gA�%�)ȝ;Xh|����qɡ�#�o2�0��s�ߗ�ົy�u�1�B"~)}�y7wWn*��E����x��:�$	
5�CK�;���#f�� �@�(�:��2�ﰫƣ�d���Yh3��Vʠ�������2�������o	ay�!���%�zSq�`�=�
� G6��:��i�h�m/�?�X�.��(gm���l������

��?���`8�����R�d��-�ģ���	���H�sJW���v+�g���-"d_�oI.%��q��~��ǧE���$�����n*Uv��
ZUT�:���4��=��m�*��Oz��,�\[P���Uڸ�&��Kv�����P=���b�n��)�E W,�tlR7L��~� ��7����qH���ۍ����ֹ:ɋ���񊊂�Q�]Y2������T�[�@`�N�]����Ǵ��J�/k�~1^4��b�|\�RC�l���r�ZLd��oɒ'!�R��w;�dx~IGT����	�hL�>�/�isLi�Z��H�^��H�?/!�-qHy�\<;W�0�`'z��t�i�f�^ܵ� Y)�Bk���է�2�����_��'o"�n:SN�(a��0 =:j��'�A���D���>E�@��K-�Dr������T�W�Й�������鏊vKq��;{"@s<dm;u��!���N`�j�.B���A*p�R4�{��5q_����:eև/������ej����i�/b��k�g�. ��g���.
��o׮Ot��\t����5g	����d�;�q�7��&vF��ϙ������x#�u��#Z2e�|�G���x�q�գR���2��%$@�-igtC�g @U�G�k�#�f�-�uk@[��+�b�<�ƪK�S�,t���<zY�� �{ּM��L`5�F�nz�	GQ���m ��y��;��?���>�7��rc�Ԙ�Qk8j[m�8���&����s�����&z9$�)�yM����a�lS@Fb�DuS��
Bw��je���et��2�h�$�mkD7Ǡ��J�U��32E1|��Cv)�VW�w۠{E�^�Wɟ��4a��5%GҗF��O9��Q����a7�7ֽ��HsGK�"+�#��T?y�v%��j�M�z��8�� �̎������V�VL��)y�G��6�G�0>�!B"�p38������:"�s~��g��{��d�7���[�+��&b���^��ȋ�6j�k@'�f
Ȥ��֥�f@��ǳ�39t�9elO���^1�l1�Pz�b�U���ە�R�A��Xm5�B���V�P�/�W����4wyiSf5�Z��&���>Y m��"�g<ȱ��ϒ�Z��0�E�0��Z�]�F ��ky�]�f���_����oSN����|/�Xκ
�O�1�/Wa�/Ví�:�)�/?�f���H�x�ө���<��ώ�E�']�
�a�6�d�	wcK���,�0�� �:��B�0�'�}��:��=�&��bS�̯4��k�!�F�sO�XnY�H���ח)��A�9�ѣ|\��$j�$���w�%�_��_��\�y�F��}��w��Z�E �U�[�9�)o@DW~F�
H�����ƴJR®/��K
u�T��˭hōp�l���A�q��&��+�M�L���A|�f�N��u��Q�=�|T�g!�p�n��Cn.C �1��EMG�qI\d���gzX���!�%�S�$�%��1j��X�
\O+"Ѫ�PX1Zˌ��.rAmL�P��2ƀ0��L>�N��a�a9FA_�!��A��m�{�*��4�N�5`Q����f��1%B+ U�d��|.h��4U��1خE��&��B|�ȳ�z�J=�:��!�vgט��
g���k�+�/ˏ�y(��ݵ��n��'S���Y�N�Ө�>V!6�[-���=�t`քtϴ����^�~.�+�o�������h�� �e��Ŏ��sorņ���$?�uv�,K���I��.�e����
����yW�j�4E�u�}߼I�}M��^.$4ވ��HN>�����Rh��ΠXl.���6��I2��l"�+���~���s�'+A;@�n���hc7�˶>���Bz������;uG��P���qƖ��7��xBy鿠�Z쒍��Ƥw�Hmj%85�F==M&���p϶Y���V�n~��j�/��5�ƌ<������k>w�`�\���"����줳2���	�1On��X\�Y��� ����DbN�F�������hN�W����\�DW�0��cP���^ࢡm���9�)�UsO��S��.F�̷��?P���U!�c�Kk�G9]
8�p�J��r��i�"�#������,s�+�E�,x�ʵ�^��ėg@|P�&5�ʐ%w�7ei���_o�M:���3������ n�<,^�do>��Lw�p�	�W-n^�r���Ѝu�).�"j;,Y ��D�$y�;Ɏ�]R/N�f�i����t�GyKS���黮����i��ϣ��(GÔ�P0��>���S �e���Z�?u8Hdk���]uC|��$��m��6���p��۳�{Ng���[-y;0�9E��O���7���j	�@�BLwJ�m�~�m����$ص��x��?bh8�(ۓ�D��Йh�NEi��cP,=$�n�5dk���F���sH��.�4?.�$�3���%=��ʷ�c/�N�	�=,��� ��T(*hV��ΐ"f`�	���5( ��	0+:�\x�0ّe��\ǣ�����8mz�\�6�EC�`���*'��2ZE�f�^��f>kV���E�)[�Rc�V�"`�@��n
���Bo�5��b+Ff~	9��� >�	lOZӈ�Ï�li>$]n�}H�i��'&մ�O�H���s��l�ˍb(um+/���c�ks�ҲbXd�@D��`�@3�³ln�}KG��w�y�� F���~�{� . ��#��r�u�R���D\���+�V��wԭ�����$j��������נQ=uf�Zx8���_��|��/y`�� Z��G�]�e0���Y�	39�&�]��?�B��*�8z��',��͢ I��p	b�1�R�f���7A�L�-���
pԕ��Be�['�
L�/��%��y��w���-O���g,B�7[��&��t��\�O��0d�'�N�譨w8&�O����812�.F��s��jNӓ݉�:8�>2߂��!��8ʍdd���TdW��-zRgD}��XK���<���X�k�%�����C#�����|r���Tj
j�f�M�M>��J��0J�X�J&����y�qe���������Pd����������yt��K��*S�	
4���գ.��4D���n��k1ȔNWc���0��0��;���1W�{�{TA��g4����x�Gm$�˅�0��D��$���ԋz38��J��Yw�;��`�78@#W�
h���/�΋��sV�\�z�ʾ^�q��5E�4�&Ϗ�\����F ����Nc� �J:�����d\�*"�E�pc�須�9�~F��Uo#��hni<���q�I!M!�t��^IhGX��z��+�Y�O//�iGG�1_�Z5c��D(�	��e%�ם6l��q�Il�;�1�['��l�/�t�i����)�3�(5�!��4��BVS/�_s�����<e��
��B~ܪ�+����玃/&�T+�+*#]���!/��a�pE@�l�D=�����&k4�ݴ��}hG]�g�%�>�e{\�DY�g��!����EV��J��lYdb��ݑ�Z�!�/�s���<Z-��MjѾ��kE7�+m��~�>� /ݩ���O5=Y,n��g>�n���4�ߩ�g3Vъ�0�z[*�K(]���[��d`��,�&�� ��K��)�
��/�:�6�bx�E����P����7��3'�,��Uoө��Qp ��^��c�+ǈ�@��٩�������� P�o�����RN�����HN�^Խ<zgD��q�=��Z���(N�۶f��DY��+}�P݃l]��#9����r��{R)a669�;�x@��$�&�����d������}�m�Jt���K\�p�]F�6�Xx�6����"lWr�R��γ9�	�Q�y�|��L��pw���eD)E�¾�-�k����w3�۳�_6��#'F�\g�@�Q�+������`K���N�S���0A�nm#��e�: ���2x8����9z���H�S���
D}0�Q�˶����.��)�$H�U�nM�6�7� ���%1{�^�9�y��Rl�#�u�+�B�<�qX���L�
�L����	�z X�WL�I#Bh-,���%!}'�N<�O�GP�@9���f�y`�ܒe��hx?`m����工5R�unj�������8�wb����W��^"4�H	g�͝ �=�+@zw�U2�>�F�7��Q湽������k�ުl���$k�{Aj��c?���P��SgZb_t�YSR 6+��:E�}aN	��}6I�d����a�o�
��2�N���N�ĵ䭼�R��?���t����x�W0:yU�b�D���B@�)�
F澚�r�Ú�cDs�aNվ�=����b����D����$�F�_{�VVi=�5h��}�0$��n@G�t�����I)����|SrGz��t��s�9d��B���N�P��p(3i9����J�DKD޹�3�l��m��`�CSnצ�@Bc+z3^��tA�������C�	v��Db��y��|�� ��a���,�(���:(W�Iʐh�ĩ�?�U�ݦ��0��U�_�$����+�x�/���:� `4�S��Ly�Xd�^��}��e���pc��$��1�����J-�>[�UenO�\�䷤}8�����k|aΐ�%h8��!�fB,$��#�r4-NlCm������O~���B/��y�{eX�n�h'�|2K�z�Lα$*�"h:�k�|��P�������u��2��9�뒡n��d�Dg��Bu���R�!��I��<Z~@H��=r�\a�7���Ce���4y&�[a����L�[T�l��>�c�+��j�EJ�A�XOɳRD��Q�Z��>��YnA��|�cph���A�آ�p��?���T�/a���}=�:��w����]��p�����o�pB{�mԐ�r2��fc#��q(^i0��
��8������5�'�6���9\�z ��Y��-��B3�� �֜��IF��9:�D(�ue��P־�Đ�q�����7���1c$�,�(�[J!��!j�7���pڃ������]�-3D����� u���$�����$�w���2�!-�+��һJ��H�-�%=�p9K;�I˘�5g��w��Ъ�>P�Wnϴ����8q����"�gkN�P�ҩA���x?� VS��zI�^Gr ���� ��&�>-��b<������\�]��7[��Lel�,f�G���
҄È�Y�M�n:d�ɅO���դbu��A�8$�$T���L�,yQ�R����)�53�ՠ��:�l��N��D��G�\m��/�<B^�9'q����5
1�!�I׹ ͽ���ѿZ�텴`�f���௼ &���:����8�
�+�t��CBx�Ɣ;��w�=��M�2��,GN��4���l�a��Ȋ��R����ad.	d{�A�~�x{���U�M�}1
"�=�eҡ�e����Y�HM&V�ӯ<�sD�s� �s{��f��k�cE����"���C��w����Yw�e��E�CB�/���~��
M�XLl"�3ޚ�O,����nH|��`�yWP�e�DBpjݡ�0�@������ؔ���XP]6��l�-<�?�!��:���a�}�Yw�b��H�UI�L�j�N-wA&�ϟΣy7�ag$-���^�A�`��Ff�]�w�ك\�4�/��z�P�	�$1�|��H�c�"**ۍ�Y� ��|��HN�����Ic�npFow�+����?���(7�1F�Ep��T��(x/��
�h�/��7�`J��u��]R@�-������WF���z)��
-�������@3�ۨ��^J]&(�����k_�ʝ��<yP���+Q��g�o��G�h���3�n��NH+o�=������tN���^!���~Z� 3�C=y)�P�n��/hᣋ�8�҄�����^E��}c�P���EA��=�Eהяo�����S�(. fb���kjM�؈��1�gzT�G׆�����f�m!n)�����˜��<��'���݉���;I�G~�(�WD��k�WI�0��ߦ'�����"s��e:&�x�2���!��=}>Y��6�s1Ԡi�ژ���f�T�F�����.P�}�=��7]����:�� ��|X�l �� ���6����( `�°��"2Fӄ����O�G�A����+������L2������\���nnT��.͸�����/$�u���
/�x��6S���\���� ��[����9B@k2�K%����#C5�Q���"����Sxo����i�F��
n�]gL�^�(yU��Z_��\��$�V=YܐP Ć2��?p�t�z4�Է�/)���xX-�XIx`֚�i�R90�%�w���ND&�ϐ�����)ڏ�x89����5���>��������h�kR
P���Ӄ���~��
�af�z%/7�).�;�i���^x���%����e)��?_s��ua)B%?�k�\ܵ�R�MUVG������{x��}�S]��fߙx��t$Q�i��	Dk
��q�8\��Gpx���\�~4TYK�&�7��P�y��z�-�+é���yDʩ/e��������m��[Yf�z��cT�kj�U���<l�� αf�������cMؙr4n�]A.:�+l����c�ʪ	M����(�܄��Kk�f�a�`K���K��*�ԟ�T���yR8�c���۔	�S�K%�LGX�P+��L��us�i{M���$W���.b��l�E����	�Х!7#x��F����F��,���	��\e�bc_!R��CY�?����/Ւ(Fԟ��5?|��a�z]<&K��IY�Q&R^����GH�$�j������R&$s���	$���k��;O��<@��ҿ�X� :��2��v��QƋ���[����l�0��[-�H"p�0�ץavn��}�����x����^��oʽG���0���6�#t_��C�S���=���0��GL��H�^㻳@�G�d��%�^����~\�z���Os��O�qoa0L�(yHX+��i��5�|�*-B�6����ƲW\�-���& ܙ�靯���㗬uS =��o��)M4
���=�d�10���e@�:y ³��&܀G��^�>��S�"�~��!V��4������;[��.�|���i��|�r- ذ�:��1�^;> �,h��㚭8t�5)Gng�RM�F����3t쒬�29�����_�nx�Ӭ����i�<�;Ѫ�[��p�x.�C���� R��J�S��Ӕ�h���7	ޚ�����*�{��2V��*a϶�'��3�X����$"w��tŦ�)ށ�`4pm�)��Ro'����`ջ	��o��M\���BM��m�t�շ��M����ֹA��;�?��b�<�NT����Jw*y"���;�t��ٯ�����*O������=f��~�&�ϦbBrg�C� @��#�0m+�����ͯV���8![h�\a��'����-4��j�,Z�4
c���O�R����O@�2�5$tV�J�|5'K�@O�f�j�ø}�ԩ��J���������,_*y�u��&mKUH�<;�#Yb�c%��X���a���:3���z94�����Ec/��
=7��?[)beV�Y��o�g�k%*����"n�0�@A箣`Xз;-��c�8�ـ*v��*Y[�*j��2�p���/c��|�<���q�������
��^q�B��A���ϕ�j��[?��>� ?�.��6�懺�ӄ)o�����[O^��.ό��SO��71a��r�_@��&����0<=�3/����5�����'=�Ez� I�9.oٓ��&��r�=����׽$����E�+F��	I��72iS(�;�6��Ҵ-f;��B�͟���e��k	z�9��,��hEx��	�J�D��u^~4s�=���|��A�'���b��t�d �wkY�i�#OV)�!�El<��?�8��4��9�$��1�+�О���j���Cy4>�<�4���A�@$��z+H6q/��/�9�-�~�m�J!|�KȈ�ړ��L/ϜҺ|�|�6�=�7o#b�9	���lw�2Eџ�w�h]�����L�)Y+��F��&�F�H��,O�Bu���"�ז��4�wM�k��B��ɵ��fZ#�A���h�/�Ȇ�^Q�Q�H.�ͼ����k�z�7��6n���p�;[V�F���y�ho�#X����������}�~%ػ��G�t��v���*i�7g�U�V���:T��ӦI��r�%*������1T+�j}Ԉ�4��4R�a��F���|Bt� ��s�#y-���)<9[P�E�_S�v�v�pJ
2�0_%�7Sg�W��޾x磠��KzF�%p��<BJ�`��;�'J^�+c��{���d�:����V01��@��Mt��+,�C9�f��mM����E��l_�2׷j��:n-!v:M�F|BD���_jo"	�Q
�(��N���PZ`��֘[�)��D+��y�,�,rj#N�~���E�`���I�ാ���"	�XX�Nk<�w�W�*�	����E0%o�V*,�b���2"����a"+���zƝ1IuYe��\6�X*�v��ܰFK�8>�O����*\��ݴL����Tօ���7�X��A0G2̷ܩ��YU�D�_���
��ݭF�Ib�V����U���M�[�l(����_̓�o�^�4	�%���ܝ�l�m��� �.`�%Bԃ�X	�"��W��p�����Y����N!GA�����<�{O�x�eÞ��9��#ƇBmAG�3��a��E����Q(�g�Av��� яG>�pt)����\mzG�\<T6�F��R� -�hX�����g�=d7l��y�y�ѵ#��7\ń����5˻�KnD�u��U��g�8&z�;�ܔ��� R^-�*��'�[S��Y6.��	�|�o;V'wm-1�B�Q��LH��<@�ڤ�/9 �Rl'���@xҡtd�qf�ց����Z}RÕ�
n�ٷ3�N��N؀�Iz��,:u� �x�*��!������X���Z3I�R�q��H�Yd�n�lS�;�r��
��A���-P�fKݠ������i���U]~�P�}�>_��'\�q0��@�v����K�V�0�ƓN�m��^��MM��d��kӢZ<�G~���)�t�y�!�&˱Pp��ß*�.�Q�/�w)�5���ݫ�##��E�H�����a��F~�܋^>�-M��n`��o��y�GJ/���A9tB��k��$�"��A�=E����fWJ�v�2|.ޠ��m�٭���^.����c����NV���f��9+����\�҄�@P#)X���?y$+���@b���u'i�P����6KJ�Y4�UQ��v�h��i[�PB��^��g���t|~��������GB�j���oVx��t�����]���]9�c߳t�����'�W�x"==S ��g�>�*�8��e��5X�aN�ǣYR��\�Ӻ�(C�s�V��.�d�����˱s��߷��������$�^�榗$����$��i�j]95��VB���Q{w�I����,1���I�#Lˈ�A����2ҥ�dЉ	����s8��r������y�a�����W]��b�af�^]������������O�"�k�c��Cv��K J��mFk���
�ua�e��Y�	fZaʀ�02p�\�>��Uq�3!;
D�]������h�.������@��&�ڴG;��8��� �j�靌��e�.ЌQ&A��0��a�X�.I@����c�*u��l`�R�)Y@
R�S���cO��]�*�dʡhU�H��lq�i0��q»ޜ{e���S����4a��Y���H��~��*Jք*>h ܋ax�~�f3τ���O�+�2�4w�^��0-�\ᱵ�J��5n#
g��ŵ���?����S<縉5;��*jꌖ�ϲ���/Lg-O�}t�����i���瀆�b�P��s�c����Fd��0�c� b ����f�0�c���d�*a��]̳'[��.�aJ��&iӮͿlH��0���	5�ۚ�K[x����0[�S����&�D�̬��L����V/{"��-�� 4Iz�<���NUfI���[���Ėtwf�8:�~Wd}�a{�(�j����h.y��b�/m�����/�I%���&T?�1���ǚQj������0槇E���?���Z_���S���2o	!M�_)ܨ���Qa��z�|[j=���
��Ǩrn#1�tp�T�tP{ɕL�Y�������Hݬ��?�<<J2M�/�E/�����$��)Cڃ��j�	�̮u@e�	�MQ.�C�A�`��_�wٛ�"B����G+�H|�P�z�kh3�I�����ޕ��;K6D��8���=3K��w��)~����Y��,X�����/�]��|�C>oP3��jd����<V'���j�GN���u*۬��h���{`!�{[DUA���6�&�=�t��C��2=exH��lհ�l����O'"|xQof�q���K�vdzS�|ea�ۧR,n��i^:A�`f����_��1m��x�o���Ь Fa7�i��ps���7����2So���y�n���)�r�ne������tu$�GU�A��N׆p�{�W�6V��.ݒ����8��?H��L����~�!>3,xfk�Ѿ{/�ct�*��8ز�˰�-�)2V��妻'�1�@3���y&�΃�`�V�������A�WÑJ��ꖟ��) ���d�^�c�j��(���P��^_��X�c�!��(r�&�]�u�>�qp)��1
%�a���W=�YlN��ؼ�Y9Le�Ǜ�^/КY��5���_�+B�)�~O��`�%���s�p�R������D�i�F�8~�ڍ�1�4�V�1���GJ��e	����'�w�b�ҽ7�d�QH׸�X�
W��6Y`-���S�x�R��p]��!�d�h��Y�bP�F�7�?noa���@o�͇�'߹9���"&Q�ӛ���%?8*��u����<j���~�	��_D[֢��He�-�3�� Ai��5�M��Xg�О4�6e?6�:]�NA��}5��F�oў���������תCBq�e�)$�b�A;���]������8H�ʩ<_j푯��Q�*�sK�V��w�}�X6)��ϒCuop v��]SK�B���v���ا�`�Ԡ{��p½}�y0t���¡v��ԠZű}���И�ON ����D��	���ws���R�M��c��Q_CH:�3x(5�$�0����\L��,?�#��zϟh\t}Sԋp!�p�� �{���d/���#EX�w�Ϯ"��e�^"�����D���K���;9�X�q�΃���ٛ߿�/�*���c��N�����v3�f��@]�BP-����}s�r4կ����� �F{�V�'�Q�	ke_e��;/`\��MfuS��%eN�]�p��[���<qٻ�`�� 4%,Z�ger	bVOd�3\�����#����y�#��R,�w֕�`��^@��A&\�^Ʈ:I���3zAD��3�߿���R�T^�;�Es
o�D`w��"^q+b�<n�!�|L��S�ج7`��K����(fY��Y�c�6פ���"���?��(�b�B�ˬ`.��!f�P�r�LVt�ftS d�[���ʎo��꘢��{J�U3U���%�]�3��z_�T�R#����/p�5=g�E7ޮk���;�����$�{@�o����axG�js�7���L��,��Bm9�tA&� P�K�?��;h؞���߇%}Q�'�{���D��CEBr���/#t����2M��`z��}���[������i{		$������|�Q����b~�aC�Y����fȰ$ߍ�
F�D����}�4�sǚǛ'28�;/�J
���g�:'����O�P,�2���y	q�Q�
�rw,��-�n����!�����*��-�'/�k��'�צ�-+�~�'1v^�v䶄.���o�p��*^b,K�����z� �>|8���L��X:�L4`��Բث#����a�����2l�[�8Mw���T9\��ݫL��uạ$~�KE~#����NfxO�����'��-`)p']�W"|(�7�!���N`����G�>�ޟ��fc��T�h��B�i�)�> F�����T�k��Z�q�9<gBE����i3w�%3�6� �X���&��Z����G�Ĉ�u��޳ù���6V�Hŷ�N�E(��1�"'_��[�x��8VA|����hQ���,��o���!��j�F��jhT�<e˂����X�r���?a[
I����f@�����%��u����� R�3,�Y� `�m6�ԔA��S��-m�B��<��j�3�Y���X�����U�P7���+�=��nB�\@��#���c
��DuZ���P�f�sM�lC�,b�
ť�R� ���R=F		;��Q�\c@��?zzo�ϖ�.�E��3�_���k@S������ ���0�^�ldz3�z�H��a��n䤷�y�n�0w�j�[䪊��SǼ����+����z��7���٧�s�L�<i��?5���(��2�VF����!�X�Q���\L�/��%ǭ���W,��d�e�2?�}�������#�alynP��2�F�L�h/�O#�|շ��E�q��� ��[��һ~��ZS"U��1ڮ�<v|��sf�	_�U�t1�[q��T�?�Hv�ld�O=�$td˜�	DѮ�ē�]w	CB����vi}��uUkٗ�h�O�d�=�J��@�&_���z��Aތ3�=��X��\�Pl��R��>uŗU}�opv�����QS3�O"c��qS`��D@����HD�}]�4�����M���@�ڮ2�U���	�=r�T0�_�����z�mWۮ�0$ɒ�i$^��2\;M�_��M.��M)�#Wz���ۍP�")G���pT��T���CE2��� ���hԡ��5P(�$�{����.Z��:�g�%o0n�4S��KgmLC�~<�F�R�O7��ru�[ݗ!W��:���j��6�DW�_�>QE(�������Or��c�cѩ��~��X�{��i�rB�#����̡��;�N_��9��H\ˊ��;���JjᲒz;D�I�.��=��/�ڣ��>�B���u-�7�(r����:�Cc�٤�����:�-͛�!�vM%Hy�"'*�V<�~@./HQ�
d��b:/F�~��͓����eC��S�����s~0u$�\P]���θZu���]��ӡ�����1��޹�V��>���Y^�/׬>����)�C�I��ol�o[�9f4D�H͓5�]����,�:(� ��)�ӯ`��W���Xt�q@C��IK��'�)jL\�yW�"����d��'��br�8Ӗ��<G�wD}KO�q%��Zz���M\��_��&\���r꿢�]hvn�L��P��?{��đ��0�pm��`
SO�5x����Z�I�,���� �V��^��w<�/P�k��e1_y��í��uMODvj$y��jڂ.��<���U�� �v�XI=���4���\� �,���	F#�P�yQ�"YDLc9�g�H�5�
�ᜄ1!N�`(�e:#�}*%��~�l�?��`mE9-r�ٟ��(+&h �����1���8��!���i����tſD��;8�4��Ҵt�X�����%ICy�E!̔�j�yx�-����B�u�U��D�&<�;Q`��Jj�	yZ#�P���
��;{2n�k'����h�/�s/�.���=E-��0��D��Ј��!�m�WVé�=�BAb�5����������։R�3�>�nװT�S��LDE"|��
6�B�l��9���iX�Bƀ�a_8|�v��灋���!JԷ�Y��:zn���I�:*p�W0��!�OLiÅ��7)3������P��\u��aAR�؆_��r6[�i3���L��/���K���#j	3�1"�۬5$���	�<FI�g���œ����	�qA�8�M�%2��ߓq�/vI<� �d��@#/������]��#��m]$��t�頞r�.`G�
���\��N_��P�����4a���eU���Q��}�ёOBl�%-kXm����6�Q��
��e2�	e�V[ tv�o�	���
d�� ��k���'O9��5d�m���>YW�v�kB\�IG¸V�T�G�O'��c6k`A86-Z���Fʌ��ͿJ�K&��S���t���b�I�9<֩Ж3�͡�ϥ��#��mT}7j2b��z���V���z���ܬ�y���Փ_��H��5�� w0�nYIg�9~���wq9$�f���O��m/���09��+,0�p����yY/sK�R��W:-	��߬�E��C�vj����,��N�7>z)�c+rg�H��3`@��+嶉T{�ŝ/����G!�FK9"�_AG��H�)9g��r���[g��"�fB�t��w��<���>c2_#���E��Z�։S���c�[�Q~� >VbN൞�W�
���e��9i@��j�k�f��u��mg95��od�\�����i)Tʚēb�N%���g�PU� ��+����y�Գ3�]߾���Xn�O'p�.�KX��i��Q�P�L/XS�����D�݈K
V��)<>ς���p4n�w����{;o�x�����O�F�/}s����W1h�2�����=;��s����>���D2�Y��.�����Lݻ6������D�cq��־��a�<Vq�<�~�����G�쬦��>ccҚ�j�{w؁�����i��i@�Ģנ=��l����k����X�ƉU] �?
�}H�d��n�Uh�}�U2ܣ`�qK�0n���.�����+æ9���$��2�3�c�=��sa�=�F1E0���$��#l��ԋ�4�~Q"nf�У�g���z��_lX�^�)+�;�,z�#�Oi�}�L�Ӄ�X�=���i�ڡY�;?���W l�"��`�"�:<�+�i�EP�� �*�r����m��}�s����z�C��(�t�b��� !�����5_ޤ[*��9>tu�#u���z�)�DO܌�6�g������W������;�8�������r=7i�����+�f�x�&��ҋ�0��u�ss�k^����^��8�[��$1���j۽���FJ0��%f��C���g>W&�w$0��$Wԙ�v��H[��e�c��1��l��+sÅ?���PO���|�z7K��xcW��z����%.�d1<Y�������Y�,l��Gu��& =�Y�w�\`���u��+I�W��z����y����	�0ͷ���W���%�*�6:��@Q�����+���mfO��SL�D�b��ԙ�D~�G�p�8��#;�ԯ�~Ӭ#A^?�R�%���*Ğ+��Dq�#�z�]ruK0�a�!hi}�l��[�-�%�ҧ !��%r�ȱ�k}y��Hd���^\� N{����t?�No��/�:-(Ip+TGh�.Z�;X������Ǡ�S6�:q�2��kT#-��ʛ]�S�JI��t܆� (P�*k��� T��U6A]��K�;?Z��o9�v/?�T�]�2k�~�VX�����t�ơ��^�}1��	
 T8ܷ]��!A�C<�`@./\�)>2���Z�ih��Lp^�����H�:�k����<��$&��� @����|OgE}���;o�޳o&�knW�d5&W��(.�y��#u��sAg�,J��ߦ����u�D�;�/�+���E�VE��)�*D����s@��P�o�x��TB���`�*��i&a�},���������2���A{���W҇�h���5����G�%/m�9F�����*X#�
t����|,<�i�Ry�6{��ZGǥ(4#�����6*	z�"����__3�N�|�\���`�N�)b�#�ݸ�}��L$l�H,h8�ÅMm�����(���:2p�4���{��וtx��6`��/����|���}�Ri�(��׵�e�\o5#�p������� `h�@K՚G���?�CE��.��Y7��'P2��2Z�"�{�"D.���)6���	����Z�ޡ��R�: �k����#�[I����f�uC,Lg �=�IE���Smi���Q��,]un�^1�Up������U���pMhχ9˼��tN�q�7����Y��zx3��%d����U����Te�c�=�.|4�D	���J�ɽz��k����Lm쳳��~R3l��G%�9���zJ�4��ja�,�Q�K�J��������$����o�;�Ni�14��^�:�Yr`��O�#5������ŻY7�}��W¶Qv
��W�e�ξ�6�@��i(�����>�!��=c��#�9ǔY)%����E<$�%���,	,�q�	�)�IG��Mx�fDS\�(pn.,��� |~B�c
0�!l�I�̙�i�T�|���?d���j]���thX���T�>��[��*��&ljc��*-5��1�����}>n~̘�1���gb�>���ip��{D��P�W%���B��<'�����k�C*�7H�cuQ�qEz)�ڵl��)5צ��0n��Ɂ5�$���8������?�I�CN=4�W��G�; #x�	�q�}g���h/7��<�@�RG�Y6{����$gns�ͣ����a��V
b6���2PF4֏��і����Hp|\��p˵���I	��i���9#Ͷ��u{���o7dC�Bsɔ�h�W[���_�#���3�|�k��Ա�ͶcR��>4�;�J��ܓ�*�M�5����RJ�dw�i���`t<�rT������ӹ�)4�[ �����X�+��7�k6b/�=��5$�>�c5��;&��'"��w=��	�L��_q@�C�8�ߵ�l�����ٽ������6]�Mm����U������M&�D������kK��8�J�D�Ǹ�� ��H��K5��P��b�FR��])�?̪�u�s|_%&%)�&~�
 �G�����ay�����@§�q�f��C�p�0r� 5���a��+����89��b�:�*9����c���8�����F�N�iM��ߤ�s�3Cf�% S��8�iTm�p�=�?!�B�����\Z˂a�J�j*+0���O��{��=�p*�/�f� �NQ�w]A|�h��­���_!��5�8m��r��G�GQ����[�-N��q�H
m�͚{wa��>�N9<�.q�U
�m�Fo�+�mЄ��w�7��>`.��>u�pJT��Z���CLώ�[?ιh��&���6�����s�π&[X&U���_��Zs.��e��G5�g��+�glϋ��<+VM�g�yJ^�u���h�����*/@�O������G>���~/X����yXf>���a�[�םg�Ł����yUW���+f�	�TS�n�ͯ!{��Z��q�� ��~�WL�NA��1��8��6X�7g�+���w��H��n��:�K�M�}uM� 6M%h�6Hg����!������hV�iX�/b%��5��Ӈ�e+(�r'����x;*��&Ƨ���̙�j;�e���_u�gscYY��3�a�Dg�A���$]����AcG��|2B�I�"�i>˺��%�e=YQ
[�K6k�p&���/�u�R/�������#�Lv/K;/a�\���C�}!<-�V��&O�2
L^�Oq�ij��K	uv�z���x�ޑ`��Ѽc �x�#�π<��'�ַ��"BF��������O� n�>��SQ�꽡=i�v��Mp%j�C���ر��]Tf��X|�Q"�d�A�r
���	��o���1 
�x6�(�6����9
"��_��u9��bx�|>�R���>T�7�~Ҵ(�7�jLM����p���L�\��餻��MJ�\@[�}���C>���;��t�Ӓ�|��v
��j�4����G[���w��]����dk[�V֩�"�ߺ��:�<0Hc7�p��P8Q�͢�6�&��U�w:�j�6_ZU���T4ۑeKMލ�9���K� DC	���u6������Z0�ٌ�Gu4�!g�QU��RP�@�D�D��VvN c#�5����{.�bx��Qu;�q����G;4�}H�U����|Jč0aq�ݻ7B'-�0�δR�c�KN�EÒ���I���c��1\��{Z5�Њ��(U�1�}��2���R���K���n���ݎ����E��c��q�.S�X��T�pԖ�V|6NOIݤ���׀rzM�P{�c�9 �����dʴ��2g��
�g�Gn ��6�Y�R^T�)�W�&�r��+y��#�Gz�G�e!��-T��G�;����N�:I��$]	��w�S�{�{�͗y��)
F���6WZ�B.��N5%��f�#f�(
q���IO��m�$�3��-:.�围!XB�x�Ȁ&K�����B[a(��]o�F*m����pHI�ޘ`�C���ؑ�6>Q{_
�UB�p��VD��\tQw����t*1xY��T!�ıb1���Գk0iN̅_�r��(f#��V�Pǅ-U$�<]!�g��C6	�w��BԲ�ǎ�Zi��x���25]�)�
�̽y��~��w=&�Ø�`?}�����
��T��H����E.K͎l��Y�c�ߒ��邚$��T0�Wy,�Ɠ��Za ̵�����'$�X���랛�r���~A���|z���4�2ֵ���T�N9��D���X]B���\�}!e���ߵ����C4�n��tN�y@�[Df[E�g8B0�j��@^a5��&���ʏ��v��W��b�[�p܀X"3r�X��q�~R�7at�0�ں�t{��n>��B\�4�"N��PI�ix޹!�������ʬ��)% �j·�w9�Ő$�IP�qY�����1KW5g�nm�*�����6ȟ�O2�Տ}.�B�le�!��S�! ޝZ7��Y3���Y�{�	�;xW6t�ļ	D�Ⴞ"6"ܺ����,�^a��f�D_�<�^�_*Fƽ�|��x��	�n[�K�I�O˄�	Q�&�^�ߨ8�b��mB���&OE�˙e���#8t���9��p�Su�C��bA���b���!��}Bꢗ�ߢ��X�]hE]�</3�Ҽ
o-��Pf>>~r�z4^.���;���;U0���`"�ct �H߸�kS�G�����M[桿Aq,ìt�.Y7�c��P>|ݞ�.�@�΀�NG�;���y>�-��
@���a��T���'��-���~���&J'��W�k"#��:G���=��wE���|_�UE7�x���|q9����c-+����R�D�<�V�H�*7�]�t]���Ob�?i��a{�->7�2挡 I؝��q[j��d(�L�85M�u:FX���o/)�tJt�DZ��`b���V�8�Q%vnb/��*T���DkN �,S�����|���b������$I�G���8>3w��*�`C$ӝEx#�߿N����:n�k�U�^��M+V�%\N@�:��h6�t�J�@!!l�3aVZ�)"0z��;'4Pt�P~l7ʯ}3Eqg�8�?o&�Z.�i���-ox;�ǁ�h߲�3<�
��-���8�&���-����J�5��<���H_-N�C�*�׷H��]X��n.��/�eʰ�LD.�8Z���&qVh񮿄�2M���$kߐ/ܖE�HHtG1��E ����bƪ��/��e��Zb"���;���j�iy���1z�ނ�]a���x����Q�*����qg�K"��P|��dR�R��y�0L�N�f�
�tòqo����6�00Sn��� N�v(f�W��:����l��C�-�5�#bW�>�q)1�gj!������z �RR��hլ�"-?ヰ���UgL�HԌ�x5���k,m���y�6�����X�Ø�w�O(��x�8B����c���K���0�ކ�w���L��΄ 3���`0��hjt�i�}�P�;yV�'R�(!���U�wԉ��2�8�>����&'�C
��٘g��r�Ul(I�`B���W�q��}����rcP:�E�sS�3��ɷ��m��l�|!ME�U�-g�|!ZI�;�z�jp�pS#S2��e��y˂��'<L
���rfd���@�"�%9n�������c*�asb�/�ʣ���H��I��"���b\�lR!Ӂ:vko�y����S���>G�}3̻��|�E�'��Bs���D�$�j���I������r�~eV{j��)n.���L!�PB7�3N����k|���
U�m��PL���a���,ڮ$r���̩��0_*"�9ضك}��,������=%4d:�=bj��7��0��	z,q>z�����L��e%V��R���8N>0�KV%��*���R6�h�Z *��`/gSEƱSՌ=&)�g�zTՔ�E��[���o�+��W��m��p곚��N�����
���?�Hz�4�� ��?�noec.��t�l����8��SRo	݌4�X.xF�n�<O%,��rg�܃[�C��
�>�T�}�M�y�ɋ��Ɛ�/.B�BXr���їR�Mu�Q�DL�GǏ���=�u��Z���nHI���V��ܶ�� �ž/��]���Ug��6���g�E�HKW��ȍ��q^�OE�?J�9_�C<t�W ����~g��h�J�#��:T�(����e)8f�kg$��*�೨/��x���r��8L6�f�ZY�iT(���c�]2x��b��*�֮��+O6&ګsj��O`�ô��Y�g9@~;�U>����R�oW>�Kk�/5^9�m0r���T�?��L���z?-S"��d
IW�FMw���C�!�Ωn[IM�8�1w��P�D]���
b�%��=��É�^�koi1sG�T�fC�Y��O�����"	r��+�ۧ|ɷ�9�rg�[g����L�܈FVtC���t�z~�\g��F���F�y�8�޲R#��j޲_Py�P�c�gv�e�����U���*��]��'1�)��yh=@�]�V�G�b�0� ��n\p�>��#�N&	�pA��N���l�t��L<���3���5vN��z��I"��iP��rh=D���8�Δ�(a6]������Qe۠�����=�;��?k0�&��#PAP\�܃mX<�4j`�e���H���1�dQ�o�l���*�G�f�:)C�y��P�9I�j��,��+ڿ��O����wc�]2��:����M3}��5Xv3��_<�6:3�.��u���4������
K�M�Gb�H�B�j��Da� D-�dR��#��q΁ 6��=�;�a��<���0�j-ނ��%�A��D�M����"���;��_<O�e��?å>�2�%�AH���>��	pÇg�:�)��P��	9�3*��:�����j�ha':�~
Iy�j��Œ(�#��H���S_�}�6���%��y9�rbm`��zO�@Kv���N¦�M����n��1����ߗT�C~蚿�V���
���.a�;G'bY�ar���&-x����HX��]:!�K�'>����׬�DZ��u�cM�.*8ED���s%��XČ|�)��՘+K�n~�0Rr-�tӱ�Q��7�� w��.��ƨs���"rd�V���~�Gn��;Č��Fz�x�\?�.^�o��k�2�.؜�o|צ�����ظ
2�w�iṒr�}����w�.�ErǶ�nI܆�~-�D5�-DDC��S�n�w�u�R1�"t���5�X���_�s�MI?���Z��r4�9e�(	r�D�7�)A�VĘR�S�g����F ��d\�����pv��Q�F�e4R�Q�J��Pѩ�����-�C�z`���;����Ӥ0(���^דZ"�-)MG{e��'���{�Ӝӝ��Cß�T��Zc��Ix�WZ���2�E;��y��1�+�ə����_�KzME�L٠�F%���<�F�)_/�̱�ꡤ����Q���h{�+X����ɶn�.h��/3�L+F̰���YY䐭��r�w��0����,����u��*���uQ��%p&n/K��jB��t�dqa-~d�<[lz)���6�A�?si�>]K�����9�
������h� B�|�:d��� =�f#�$�V/]��
�<�ݮ��K Ȣ��F�q�g���)\jN0�����,.��R��!� ���fR:�InJ�$81�_KӾ�}���qP����Hn'�^-ܣ"
��m��!���ӕ���Ӿ���T [��?�Rx��sw�����6�6c���$b��?�_�����7R*��e�%(N8�4�M�X�6�0�_��O�NL-��Ҽ��QZo\��/p��hCټ�(�D oO�e3�P[k��b�:���]�P��N}��9�Ӑ�]4:{ȡ\�e����MaSm-�&j ��~*g�&�K��Q�,�c�D���s�F����Y:��T\C+f�3���8��]soR�����JMWg�\Ic9����[���0a��@V�7�l��9[��u���3MΔY�$�@"%��U�b{����/0w��%���$�d\ �|86*��5O?�)��Q�5Ԁ*��:�Tq��2Q��1���VE(���O�V�_d<Nv�Ou_OI��-i��W��є�U��1w.��c��5�f���<eǽ�Ő)ba5J�4T�89ꃫ_q��9����^W����{�����|V��W2�]Ν[3�g��� �t���s��}Yb�~�/�ãl��?�[d8-�=��{]�<��ݑN���'߂`Gŝ�z��	ΌEu�g��Y�� ���7�=�^4�֮�	;�OȖɈ�k%��1�W�&�˥ć�9?�-���Y�'&[]�ܺZܐ�N(H���n�9H�S��)�zݭ�
�>���df2Wb�ٿ��' (�D��T��8���C���p�;��=@7���A����85�ꉍ�%�b�?Ƒ���`?�S4�f�x��+9?�z}v�����*Zx���]�$�0A�u�9�����s�:L6�ׁW�1�dh���. ��%��Yh�P�xV�y*yH��� ��_��t��U7�TA^��XD/>�Ci��#����fB�Fů���}D\��OW'��?�{���cB��'r�����/�����tr��*O��w��7� 7�f�M.U�qy�F�G��E.�����
d$^�c��<�q�1Ș�����}������VR$ż����G梆@dI�P>����U��X�*]��W�p4Veܛ��'�J�:�����b�q�/����\�3��s���i���!��Q�1��$�4���c.���L�H�%-5[�z^'#���rɛ��g�	g�hl\�{��4���>t|���> Nq[w�V�h��'Z�3��~B���ƅ����u�ߘ�(A;�$������.��x�eH��b���\4����Ud�ak��^0Cʪ��~Q:�����K9���LL�pL���Q!ϯ�E���U
��/�e��C���Ȧ ��FB{C�f��:R���g��7�ST���Mʎ�u��d��j|i�A�i
5 �<j�B��?���f�Q�j��zA֢�|��\́4�j���c"�7Vh�1��2�@@�7'@|�v�*϶ =�����%��I>�]���w���S�X8N�-�yx2sI43�[b{3��^��0e�Bw�c��]�����(�YϞ�e�g����A�8	��
L�cgp瘠��k��������s��5Kc�H��Q?���|���-&��㶪���P�K���Dj{F�Z�+��J��Xe�n���t�f��(�ZT�#�>� ��B� �6闳Ԝ�����d�(�2�ޙKR�e�d`��}�e�(0�'���]����D���?3e�np`ʰ��Rq���q�QR�s��}VC9�����j��1���~]Զ�4�M�}0�Ic]NC�"C4o G�˂Ȑ&�ìɿg�\V,D��J���u ��Q*����/����������� :΃���5v4r�ꏓM�Z���9���l?�L��|��-UaD
[2�U^����|x�e�^5ɫb�{�P��1�
2��3bF|mD�G1���)�"��A=�+ٛ�|#���1~oE���<r����lW�1� ?zD�}�5���\�O��l��5��
�J�s��Sx�ه\Z�U��L�!�:�^��|� ?�#^q}C'�X��I�"8��%��(j����M:�<��cs�v�s���0��+I�9P1�o��9�*M��D�s�����{�mQ��0���,N��L�)o��	
��m�n��`����L�}|�(S�0�Y}'pj��&��FT�'���L�����V�-kfS�����I�x�s�N�,8#��j�dF�*��SN��0�t򒦁��Y<���mg�O-��9:��%��@S���уw��!9 J�@M��V��������l[�y3�J)��eoA�7�@��}Ȍ ��b�|I},b/��̵VY��tQ���)�������\|�D��A��P6��Rds5���0e�ҕ ��D�m��Ib���Ѷ8�\��Qb�<*�(��ˈ/�!����uW�[��Ė��E��2 9�RqƤ��'�C���Ք��[�P
>�w��u����܀��.#
��~N[�w6{��&�Q3Me�uLXxʋ�w��zX
��!����.XHFu��4��Ƈ��i����އ��l�l�aW�,U~L���J��m=Ӯ���l�h�Vр���D� �*�o���O�G�w��J�3���8���WĻ�)���@	Ŗq"'+�M����t_ޟJ|QN##%'���4�������U����ie����U�/��_9�_�{(F�'ʡ.��1C�p�D1�"�(��Fl�e4%�LR]�9�AO�B6I�u�a�Wd/�4����Y��./S?8^�ʭ
��f���/���Zvu�+���9��ڱ��;�"A�h���(�yf��$��	E��5H�u��ҥ�	�!�9�����PD�,�Q�ޑ�k��)t��l�¼�)4��tx{����Tʄ�j� a�6O�$��^\�;T.Тn��=ǣ��������fR����	�QuY[2L�v磔`��&w�ڝ@(v�r2ھ�bd"B@�ZL��p;�'-��0�8 ݨ���22�4`cT�K\7au��2�D[1���1�b��e�*��Nwk�@(dO��P
��U���Bwx��W�����jz��K��4�P�g8]P���Dn��[l=.!��ןS���
b�{��6Y�"�q���K�����umH����F]���7j�Yrq��a�v�Z��͔7����Βm@0	Њ������w6U �{����a�2?]E�_j��Z\�lIXV ����Q垷����G�9J��zp����h��Eƚ�je�����O^��)V8lᑐ�P�y:Ѳ[��� k�X|�gP#f��x4�$���q�:K�5(��jnߍ{,�R�G��0�ZV]��G^��B󅿡�up�pF;]7Ȉ��w��w�����)�3�c;tS�rf>�XU~+)I�$_[��~e�aہ�q��@P{w|�ى������"H/�Ͷ��wIO{��E��l~=�4ܿ�"q�e���Q
cO�d�fQ9��ʛA��ԗlŠ����v�a��d�����T}����bbF�ȉ%�e�+�ٯ�x���#���h�˗������T5��>޹^�>Y*H��v�o�Q{_��3v��k>�m��)Y?d����t�C���c��J��m�v��ѵ�C���c&�����N�����O6ɋ��*������m]*������!e�����:U��z�w@�|E��;ߟI�����b_�럠�>��ʐ�z}��CS�e �7��<s�u�H��$7��-`D3�����8Z!�?��i�G���  �\5"
�*��'�y�����m���[�	C3p0��3I��@�0a%)�b�tYQfk��H�%&2)�X���ݮ@�C�S[цldLQcl�sٙ���fW��U��p�]���0d��	��G�Q�X�s�K�G0�z۴Bg���;��?�N���Si��X8=��m�e��}��ϼ��,F�nɹ~v���������/ЇӣLF��!6W*Ӆ���is�fE�λ���6��qBC��`AZ9}K�3��EzP�_�b?��#2�c깥+K��;����M�Z6;)	� �{��T�^����)�ᡠ��� '.d�"-��y��w_E?�+������j*���G���R��X�Ҋ�#���7�e�w��p��M6ۗ�G����d8��!A������b�g_{�xl��*mW1#���*�]�]��q��Z�Ri�����5���>|���ɤ���t[��?��t�Dxg�8�)<���B�w�B��dK�/�w��C�K�ĥԵg���� ��������{�a+@��j6�����6�~���4*.���u�R�t�1ch�OY\ �"[j��j�ox݋@ٝئiA�S���Y;"�	7���S>��Z�4$��	�D�[j,�ۀ��Ë��؂��t/b�Г2%���#�f�����H�ib��v���и�`� �;��j��������+�0tߓ�>�����3wْ�N��r3zPm�/v�(���~����T�f�ܥg�2���5���i�nZ�駈�p#z\5 e�0{~XH!Z%��d�m�[��j����1-�%��v�5%�A@������\`Pg"M ��<���N���g8Js׵�cѫ&�Cրh�(��pN�k��ON�m�
��<��n�?��KT!��y�4ڀ(��R5��ʮ�ݎa��U>[��T$B��_7&7�٪u��
"�&��׷���8oi"3�<�ii��@��+�C�#�ʾ|"�G^�2R����8�=������!�~�[A*���I�Jv���_Z#?s��(6��5����ܙP��:�DUUO�1�����x~�! |Ť��qҔ��`O_��TT'B$A�=kY=U��#�-@����<�Q��D�p��ѴL�/�}4D��
��n����Г�h��k_0HF��K��T�+0nK\�gq�n�I;�[:k�6(r��zp�mGrJ�b����������6G���z�S�n`��Jɓ�6Z�߱A��Fa�ᙛ��咿APĂ�Ŗw�GV��>�`�]Z�ɾT����������r8��n4V��[��,{oc� ���܈�ظP�!Qf����ü[xFY<�.��n�.�۹��K��60&����Z���j��d\Mo��p��;�����P�s�P���g�Z�dX �u�aS����O�?�_�QJU�Q����;^e�V���127vJ��6�����)nf��d{)T�B��RB�%zX�ٹ�,l�����g�;38HFy�j��+�y>�(��U@��m�����#�U8��_�!�pO�>�������C1���J�-\=�U���j�wa=ǻ�)�o���vG`fiا�$�Y'�\�G2r�5��J���h��K&q��v&D�rL���V5F��7=^WX�-�7wߧN^��8� �ߍc�q�s�!���`SX���f��U�:�%��'�P]=;�`?���M�fR)c?5����7��3�2?�Y �>5|*�kg<�X�!�4`�h��P�P��ж�$R���lL��a��*M(݈�
�����s�i�
_��GvYڵ2���5�Oo�����ܥ��d+��w3F��Ћ��X⭜�
Xj�mj��DO�C����:c+ƥ��Q�WRE;��"��W��n$�}i1��j}K�]Κ��:=�8A*7єz�QԹ�5��~U�1��fA�׺�����]�e�pl�LCw�N����>4�$:P�7�'�L����@r�|��ջ`�M0ј���	q̑�<iqk�cv�f�
�8�g8�u�f��p=��g@�+`��F��L�o`����!�~Rnv����+��71h�/ ��S�1�U�;�)��� ������H�H/~� �NRq|�֯�<�+���:��x���A-?dA'�O�=���Csdx+aX_�B�Cl�&�:x����%�Z��M�-����*�:܏!��c^��Y�]�����Uȃg��I�p����&��d�n�@9�{ሧ�:�XZNO�7�j���f���՝�=@�jHD��Ao�C�hL�a��k*}ZD!�L�~�(�{�x��`{�1�;�	8tƉ.Q���'��'���_�ҭ�0�oc�D�"T�ޭ��'x;� u���G:~�$�s^��oD%l2�	U�jP�AJ*�;����?3d�v��!���k{-]�׋����TCsM�"ӽ�ez�hȩp��'���],���q���ؙؓ.�q��a�<m�'�[/O��C������DE� �ɠM!B��\Я�A��2*�<�utg��UI���or�D9��\c����r���	D���a��V��.#9-�Vt���i�F�\@t��Q��A�Q�� N3\=J���Hm+yK�����gF`�Xw�va=�I� 5�~�Ƚ����V'O� '�Ln!.��0���׮�/y�KQC@�~���*�U�\x�77b<�C��@��&��X��)p˦��=�vBlf��a��bS�;0����/����7��j4H�q�)]yp2Z��dG��r�Ѷuq���+ۥJ�0V  P�$!@Ъb�
'K��d�)f���b�Z�ƭ�X���v��{τ\R⯅�H����.h���yRX]i�?!�np�c����^t>��愂}�:oynyE%ȭn<��ܕI�jH� v�l{+qCIi8�L��u�{<�êyY����R���-<�lэ����б#�������0���FjzZ&��}Ń�bJx�ku�D�܀	�^k�.P�D�sE�X෉���z�������h�,:��HN�w5�o��#U�?C{G��)�^�qB�)�*vޛ7�1!�mǢ:_����6'��NЫs(���~.g¦�ǐ,ySc���)�!͉�(q�r�OXǧMc(8��ɊU���[q��g�������sG�c�� n�>�%E�տs�N�6�Z��HΙs�>:n���T��ۄk��JE�05 zqD�l�h%�3�J���Bm��� ��*�S�۫r6yپ_W�����M��?�\۾�å%��Fh��/ޜZ;$q���լ#6XT��5��O�n���O�_��}�If6Kr̯��Q��`�=��ع�6Om��r�����j��7d��~'d��ѵh��Q̖3��sv�Ձ���0n���=.��;�M��j"p�hF`ʂ��H`������[��z����5�#�Ԓ+Ǿ(5/�l� �չ��J���3���b���o�j�2��������`.y��Z�� �o�!�Ft�v
Ϯ+�c�+�B�Pc~��U���9�,�\w�ǇbQu8]��:!��f\>�9�Yp�C�8�ؽ�L&W�j�57��XA���4�mp�&�A- �ি;ɨ!��T<`�gMP_������@�Є�����&T�!?5�I�A�X��LҩK���D��i��H���5�
��՞�-[3߫l���z�#�J�d��=�j8��$��Iܠ!��}�G �����C���Dta ���v,}��|7]���VX�P�z~iTs3�#s�1��� <}�����r�7I���كL���_����K�%Bl%�H�LgS��zj��3���ݳF���Iȧ>���1��"Hv]7O��vjJ�5�B���cx�yJ���/gwVvs�E��������*���X���%5�x���·�\��n��i�ٖ�\���qbOz+Q��n[����\t��%����l��u�Ů��;��x����JH��wOD��Zú��[^2*JKy�%
P�k{|��˖ ��P�]j��֗�m)�.��uzO����We�`�Q�	d뉷� Y�e�P���TmK�rF+\E�� ��B�p�[|��4�a�郥|�"�]H�GIY����o6f	��˳f6� '�K�h���� �~�xXe@FH"e�i�$�71=�O����2�v�PWXꀱ��&��L`sx[��2};����s�i�_��q*�9㵬y���t����ˇc-
�
qQSPhSZk�����ʅ�b��B+P<�Tzd��b�نj��G�?�x9hϱ,-�O��?��:�,Y�V�5��ȩ�	���d~���m���9R��pK����f�Hn/���1^�}�)���Ǻ8�]��㵹9R�;mw4�g+'��=>��cЫ��y���S�[D��)�b��e�]�f-+f�&4�_8nT����uN/�rU��@������'��0;p+b~8N��8����X�0WW$�`vL�Z�C��l�ɥ�	24ɯV6��:�׍y�����>���:"%4A)}Pݞb�_E�9^`�s�$������Nm��|����8�UA(��,�	�~����b�|a �Z&��
$�b"�O��u�Em��1��I���mhʗ�U㽑͇!}{��K MF�*.�
~��>N��W��~~���3�e�@��$;0Ȟ���xHݯڅ����H��'P�S�#�`1A�_��Ѡ��5TW�tw&F��~b�@���S��0X���e"�cn�|�)��RoOZ�Jڈ��U=~�Z���q6H�U��J y��6���ˁ@̝��:S/�6N��{�]�8�P�� �ǌ���\FS~�cv��Ű�;�{��e~�1z��Lp�����G~`_�WO����?��BM�����b��D��sW�gv�D�o����v�����)T�{�ܱ/ӝ/}�z�4�_���/�a�j}cgi�}WD���r�ff>W�����-0uҹ�Ǔh�����d�d�!К��./Y�i��76ݛP��|\�;K�2��g�����Z=�*#V� 7���VP]��
���+��v��c�Sw�@y�~����@K҈�Z���Q-��|���m��
�z���!J�;��4���Ǿ����<�4ҹ���Z���w,�
��ʩ����1�f�:�����B��|�^���dG��T+ӌp�_���L�mf�3�h��ra�����&��T���� �b�H�t�ڜ5�D��.N{%�w,����������	g;�$�!F+��5l��Q_��i�n�\W��y�t�ab�`��h�i�㑷�ԹF��/�D|������5��H(:�	΂�%��ReË=薫�a��T�9���a
��o��@�dR �eO�:�7Y�.6��� V)���2����E�n}?@��/f�8a����-1u5�9h�?���vTiYJR�?�d�id��$����"XJX��d{8�h`�V�x�or�)�s-��J�nP�&ݮ�w������B[E�#���/��2�!]�I�\W�FFT)��s���R��|;�(2��q��w�L�]�oy?o_���lJ^n����L0���`|Q�� LEǀ	�p�~ܟ����HvP;2�⍡��\���K��Ƨ�U^�:b���Խ�����Bj�|6+�ĭ#۟\���)M����Z],���xlf0A�!�U�ѐc���S��{���J"���3��2v���<�[��mOĸ���✧H:n��g����hّ�f��T�E|j����������d[�������Z���Y˧��
�ҏ҅�mo���Ճ'���:��QA8]�Og�Y4ų��M�!=<4ȟ��Q&���ò<l\f뢝�;��ӥC�{ �58bao���0@<z�$o��=*�1����^]�� ���Gv�&n%d~[�\蜋����rs�(��7�/ܘo��o+8ڟ�шg!(�  ���,���#����ڙTn=La���F|}�y�Q�L���V���*
1Q�0Y���,����@�A���D-hs�8�:g�����ܡϢ���&d�ӣ%%�j+�!�`IF����dػ)���U$րZt�i�A1�=�~ؿ�F> t�Xyv��5Nt����WH9,�T%��YD�>8�YSZ�A�#"c~KO��Q��|�^_;7\� Fv�\�މ�u_�7��:˘7�{�YvUH{�9�<�w,3G�
d�O̗<�!��43��14�Ӂ�K��ť_�,� T�(���!3w��$I��1Y���U�c����mH��^8���<���0�	sRX�zK[���l��`.����P������oR�2��\z���jZ���W�V�����E7��I#J�A�@g�}�e.�$��;�=�Wʔ]ȃ'��A���7��y��
��z����x6M,]�����c�k�A�^�7m�'-���(AĂԪ���l(h��k��+wM;[�V���+�]�D��Q뤚���<�2�P��mW��k�5�3-����/�5?��/eUο���!:T�����k6��,i��NP���3
�3)��b�?Vw�|����ܮl�a"��G?�����B��-�.^�ֻ��n�V�yծ�y��{�� 2p͎H�ȳ{�G̲���9Sm@x��ӑ��zB�<�_�Q�8��vJׁ$u���CYF� ;�#���5�.T�է*�fX]X�VIE;6�,\ιO�
�3Ш ��{Y;ȟ�����&���IY���K�C�q�+�3�x��/���Z6ؚ�U��m�X;�w�-���x ��F��J	����4b�R�[�%���K�~�ًN�;H�dc�/��M���A@R��	���U-�H*:����2J��G�c,�u��n�b��7=�:H�jYJU��+��=L�;���-�'�o �;�Q�M�Q�αg����˩�{&���I�Fjr�B�<�t#΄AQT|{rRz4п�S������"G���^��"��qa���-�<�y�:<�S	NJ�/X��4�^�Ap�Ӓ�!�%eH���7my>�f3�Z&+��� �����ŋRY[��S�����!T�Ŷ� 
m�?���p�����|�}}1�_*�;O|�4��律Y�mb�9�Hio�c��_O�o�����q���{md�"2��5ڟЎ�>���AJ�����]�^��"�P�DΑ��{K�m����x����`�Sc,u����_�(S�W�d� �܆�F�4����������5#1Z�tԧ�S��ҵqı��&�'y�e�y�����H���wv��2��YC�%BC~���Z`�ݗc �Pվƚ����F��t9搜��M��Py bMY_����G�7����0 �)��l({U.���} U�O�#PԾ��������z�|21��	P���w3�Tg�"^'��Ffd�T	ۄ�f\��MQ���=O�*;��VVh�&��Ӽ.��1zzd�~��ȷ<�qN'�PNv�|RYZ�
�E='#oJ'9I�n���'���͆�|�3�#g:K)�
[�])���Đ\�H\'k���[����?�v���2��V�F��bm�9Ή�jCF:I�����]���i�LKV��]�<�����Q�"7��v!VܞQ{
_A���cy�O&�0ɖ{�v�6���v�����
�\�b؈�D]s�t��Kԕ`v[�u��z@�!�a#�@p�O�&`��ֽQ]�\��]��<>��[��9pI<Iu(�}���J��וng���E*�N�[{��i�Ӌ[�)�{��JK��zFMgpLxST����T#>��~A��Y2��:M��	��� �����U�4��F�D��!��z�	�PWf�y�6aW"l��M<�4j�;=D#mp���)1�}��Nk#<�f竌 �|�6Y�	� 6:㈈�HX�����1'������ `khj�
�%46�����O��1
دQY1�(�'�M!8�|���K�1� 7Z[x���{�|�K�b����֦�'nO��>�e���o�l$��߻��椶X�)4L���;���L�-�z�$��-O\�u���l�NX�"}�{��	v;�bv��I2���e�XylGZα�s��X<A>�$
u�?�u=#n��v.�CF�Ӏ}�TU�gH�A ���!�W��a�����w�<4J��f�n={{�P���Jdd�BN�+4mk���v�L����,������?���9�x�x�P����*���f�77�`���i�t�D�F����"����#èA=��I+<t��f v_��I��eqU�y�+�=D���`l��Y�����
GL��[|r���ɭ��"b9��T"�X��7�Ec@�����?T�77�8�OQ#�_�Ta�a��%��}X�`��:�bַ�:>�K_�eͧ��O��O&�>U"ц��;짅����;�H��`��"c�/�']��|f�W��/���\Z@�ϫ��Y������eA3�X��`�`ay��@�c#���(��srI�g�'�g ��ʫ6�Yrsݞ�3ŕ/T�,�V��A�� $��n�vM�0�P�}�����f� E�
\@
MJw/��/>�k<K�N��G��c��dL�M|1�1�ž��ŏ^�����~�ig�7{Kф����FEV�Ź��`�y���Tx���C�~L��y��|�I�$~��w�=*����[�:pf|�[�#9��ؿ��o	�
8ln�N����Ȥ��L�����2�f_�����:� fk�\&Y���i�M��Ʋ���媼���w����2�]���H�`��8��Nelbr�:p!ƽ��s�C�`��]Y �����[z���8�Vm��W/��J��.3����+����]��KP՗�r?9|���⹎qͮ�v��BA�-(m�I^�������5�f�6���|FM���(P`F%x�_>�� un��2�)�'�W��^�F���)R�_X�I���s.�%���D,:���j��~�W���j����1���p�yβʬ>����0�ù��·�W^7i:�v^rm���I��0����qS��Ʃ"W�=�צK�D',R��1V�E��1�5k	B=���JCǇJ%��z.f�����ׄ3'{�u����_�wy�1�N�S	�6]����I�YK�@$�a�U��˅��)fq��"k}9JAp(��3l_�L�	���������`	��T�tz�Kq"����]�7�B�g�:�[��w����_9�aM-@\��0w6"�%4��c��i�]S�A�\կ��w�c+�I�[�̝�䉜�UI�\��U�L���$�Hz8h\) /A]3��G#� ��-�e�1�L��,��K�-Ŕu/���wО���ޭ���&�s�R��M�����	<�ž!�j�����.*�>
1��]���[le���ƅr�9�c?�C��է�SH;(��1�1��\��L6,��^�`��?�-Zg:�ߘrBs'W;秇�ˌ��ݖ¨OӐx���] ��|fb��a��wXc>ޅ�a�N�3���c��6�l呜���ܙ��2��������R���hWܛV�5
l�4�o�}_�'�!=���Ȑz)�%�����z������6Y){C�Md�%%4�8m��}R3Rk�ҘVllL=�\�~0�EO��'�P�E�f�Lj�>R�;NXn8k���p�7ߕ��+t`���[�f�*�1�67���6UĀ�ݴ��M�8R�[�YP���Ɛ1�
X	��R������Zh�!9�e��/������Pq�q;�RE���A�r�*鉧C���?��wk}����qpi`Il�IػY9c����ĺ�3��g�㓅���̦V��Z�k'x_���.&Q����H@o���ӵ
'�6X�.���>򪳠>�菭4>����=����)TL��p۩� �aLbT5(�Ψ;)�m�}v_�R��cP�=~
�na�U��)F�n���=#�s���������7�Hc[�=��&��=�w��L�2��>��1LD�xtg*�SH
%�\.�_���3�-,zߵ؟
Ԛ�.���*�@d����g��r�%e�>���Ƒ��2��tp��K[��mp�j�p��(�Eu�A��Xb(�DP�7�����ގ�7���+�Z���)�]'+�A�<X*�B�	�3H��)�~FI2��
��um�R�sf}N��df���S�����\�J��"�c�&/t{��5Нu�󓛨����L=]��C���	��}f��D�Ʌ������BO�;{^S��ܒg�ɜ�Ev@S"����hV@#7yA|�%S"�\�Ӏ���E=9��Rs�y1{t���)0��_�y��<s�m��J_����4֟A��:�`�a��lO �D���#X�lwqO)&;�H��pӟ
C�H�Y,^q�����8l?:]��$�� �d�\�T���&1��׋�����Ҍ]�d@,��6Ŝ��x�W��BW/���b/B��n��x=/��|w���$���ꎞ�GP#�� M���D��4��ˌ(�"�[�^X�9)nw�|�-G�%�D�7�,뫦uS�+dnE^g�a)��������X��K�z�G0�HW�YȽ $͇Z.�M�.�G>����L��~�A��2��`[�u���Mq���	2���|��/��o��h~�N���t�����x�DqB�k/ F�;���C̜� ����)z"ړ���s"�)Ȼ!��H�¾ى[5��������Z(�\�������?�{����y�@[Y�Qccnc�ۥƯ�lt�*/R�5�|�u	��fo���<�{��U'?}q`�V�h��[I�-D�f�Q`�_�E[�$���z]�����D�wXn�%�'n��LD��d����ג���{�����~�mO8��Tya�~���vP.7����Y�G�%m���Zq�/U#>o�X3�<EW!wg5U �PEs����9b�R�R�Uk]�Sѱ��-"����5�J�*�pQ�y-/�RL�-�'S��7�1�I.FR��T�b_Z�Y}����N �*��p�⹦ �H��r�}�Bu� ��fA���~Q��=嚈G����a�h����~�\��~�Kz��2j0��G�-[�@ �'�hl;�����8���u�䞟ȥ§LO��-�[�d�y)^�v.���s�Ԏ��(�ǭ2g�#9�d{�&t����4�4B+����{`6��H�K���a9�����"S��[M�rW"0�?~�NL�e�{�eh�.���7#���	��}Agb>*�i��𦙒�����K�U�����y̸�O}�`.jK+t`�� f���o�,+L0�r
�J÷�P\�!���k�J�
�	t\y`�D_�Ql��WE�X�a���}q�b�WFAO x3��cٙ�kt�������<I���0<�΁�)'[g����kH���!?2���K��w/�IW��q��)+I�y�+���:����3��'�?������$�U�Y$GZs�1�=K4�2�2_1�ݗو�Ī x��Gn�0���lkV�?�U�%Hàf�AWX�d�Aш�׮�S�s�;��P�Y����� Ym'F�-�K���0�N�\�t;�V(c�r[��>f�E7�F��<���ᐙ�M8`�8��N;���@X�����O�%&����r��u���gS�����$�	��=Y+�)�(��(��p�c*��N����=������F��K�o/��魯�Z3t����&pR:Ux��4��}���Z��	.d��II*��
�v�u?zM̃��r�"'/>\�k�����#�$F�Lg��Y��^�J���3<ҵ]O-�;�+�θ�|�;	�|��RQ#��榭؏��B ����}�b[�b�1�1��i,�1�qrfq�td���_@���eת&��h��D(M�5������T��z�7��t_䯌� ��9���|Hs�{�A�'\+=��7g�h�����.�P��Ԟ� M=BGp�ޔ��=@]�g�v�)�۶�MB9�S���0��8���RκhW���<��}���s��́>��z0��\�|+�\�⋷S���z�`H��,�2�a�U')pD?���ěu{�s̛0K��� ���T�8�Ri!lE0�Yr�-d�$��O��;�M�6�f'S�VYr�����ե�L��%���\ل׉��.�����R�4%8Il�����������%��+.���F>����kI��6t8]�B��w%���+#��4�U�y*��`�
�fn;������k���̛'@��c�'����.����@ X��y��V�Goi����<��Y=��gIm�Po��x�q�[v3�T���� Djh:n�+���=Z�.Or!-S���B,Z�<ĂY��Z#��J-
���#�ɣ�ƶm�uT������b�#����C[ʋ�/I�UM��3��qk�I4�s�+*����uf�_�V�l%�7�]�͛j� ?�ПZ��F�AHL�oSKwݺ%�.��{kB[��)�����2ouZ�[Sok�e��Cl ��%pߌ���!g[,㓽H:F���^^�	n�.��_��=v8�#��X~9�j�	푸2x��(�a�
4:�'�L�+쉦�IEB}��{��J��Ɛ,��?#��������r<���2��)wl�w��٬u
o|�׼�2I���;ܾ&x+�݇5����t�͈s��BM��J�Qp��^ť҈�tf^��3�h	}��H֚�Nl$��1�rJeo�y�F��K�����-�$'f�^Id�]��۬r�G�Saf�|�M����r]���2n��z��$O�h2�׵λ�nzU��ߕ���.�[H�W]Gd�\yH�T��9��1�B��~wl&.��)X��C��q?~aWUw~R�=1]���-�W��o��z�h�:T���~PV=���'��2 ���oz#��<B ��,�C�k�*���R�Yy��cb����U��Jh֤b������W�ym2�e ��W0��z?��'Xe��n�=�}Qm���<���u�N���lR^�>^�`��q};��9M_�l)E��]�a��ӱ�L�����ɟ"N��Z��]�j+���G	��F�[r;�u2|�nc��ٓS��ïUz�sk����E��ez$t��`�{y�Kh�[e����wDeL������C����`�r���Y&_r�;�rW#�f嵹�Ofм���0"-��"]�N��MZY������6f`�\��8PQ�v���,\�@A�mBt;1+0ɺs䢰�	W��!�X)ɷ'���ׂ��r�DR�Öč��.��x���� ː���($s��CO9�U4_��`+��^�i��(:�T6�R`.+����� 鼱�T����k,I������ ���t3�G�jF�T�z�N��jM!�&�>��	fV��/�y����/T��s�ަ$[5����]6nBSZ.l�	�7Q�S�;��$^~�w�d
73�q�9\�i���Լ�v}M$B�#��kF������
o��H.�jdN�rK�������|ܠ}��E~�n��	�A�"u�lt�QVj�N�4�'+��[����$3m��
#�O�;K�6�+FF�<�Y�	��K0$0|���T�����+y�$F�S�F�Ȣh�i�P�ռI)�܃U~Ru*���f~=���Vl#+���&J��ky�wp��8��ƽM�چb��5���U��;?@��2v����(�΁��T�ɋ��+gL��Bz���t���n��4�Z��mH�)��Z��z�bhB�s�>�_m�+��C3���Q?J(�/د�S�����9�B��oo/d�E�LNz�K{�FhJ�A_B�3��nX��'؎W����;�j�-F8��(%����M�uT�E:G��.�x�9q�4p����"�����i+(�Ž��_�C���/��I&9��+
���~ �m�M_X�{����	~}e��I� ��b=��Q�B
�� ���L�k�s.�C�MK`YN�a0�&;V圹��H��ZOG��+�V����r����HM���L�ǈ�-�#�� (���@��X�4�W9�(n��%���^<������2$?p�n�}01}�����"C�yVO �"e@�ҿ��
`8�t�)��S�ԖP�~[�[MF��mJ}���&t�s�OuN���D>�5 �i�|[3E��I��bז�A,G��̿!G�8��A5���c{���86�_!<@Q~o���.�[܏�S �Yx��R�]���J#�<��DK|�S����ou� Ԋb��X�w�����L~C8�6��c]J8P{�G}$ٮ�O1@��$#	+f��F| k�����<�@��E��9@��$��*������Z/(]f�>MQ/���ʊ��]�%>����o1�7v~�]2��2�=K���%����yi�������k���1�8��
�)�wg�'�20�� y�Z<�!3~,��"����qw
�� �����
�ݷ%����:���dud��]6`�W��Q�Ì_.LL<3��ƄN����91��U@�.�H�9��Ko�ɮ�c�.�)L)����rw���,��\���o#�m^�ߊZ��K�U��;#��p(�+���d���[�G��-�At�N᠁"��͛��Jb����f�����'s�s���F`�5���R�NOX�w�C�&�M�9=j��ш��O���uT��^[?r�p��랫H�T��T�ESD ���(�ɢж<εj��pz�Qn)r�^Zp#=OG���o?v#�H�37��6��ͧC��q$�)�P�7��s�<5k���-���yX��ǅ�W�ం�$�t��0|���`Ĥ-2�[;�����@�.�P @Z����~3���U�Ǡ^N�!;�hlip]�>�}�u�d���^F����� ���:v�rbs2ʠqE3L�?j2v��ˊA��o�HK��VΈU�`� ��'�:^�g�D$"�Om����I��q��0����q5f���p0u��h˓(xm��x!5�����L�����<Ngo���0A�HL���%;�D�x��4g�R@-h��N3����J,�ڄ"���V{�X�A;	o�ҰGM���4�(�H�k�@��"z�`��c�[3_m�a'�ef��K$\�:ˉ=]gԥ�[�H�]$@���}�À"MG��^�C�g�<t���gw�<�p����9ߢT�χ�ě���nc��Q~@։^�gD�����)�$zEf`#|�,d�kΌ(���@��Y�E��E_��8�J��ۧ/�܆	C=��7�����`�l��=�pcU,m�M�����nەX?o�ƘZ=�V��������/7��cxQ杜����V&� �ؖ������5�Ob���Ȕ�[:3�az�	B-(Ɲf�k?�����(��i�/6�=�i[ݧ��:�>,M"�ʍ������d'R��Wg8� 5
�c�`��>?!l? 9��H�d9NC����6��4�ŽOAB�$���-4P��g�B�.Y� y$��9�o`��.�'�<��
��=������k�"G����&���B���ru�m�{����I)Np�l&�"jtw���dj+}8��3�\
"y�������G���u�g}6��u�`�@))߬b �s��+�ݯ��t� ���'	��	��'qɾN��.˚̶h��i>~�C�T�.e��#t����^f���Y,xaH}Ȅ�lߋ�ԯ�q��_O9��Hl���̹ƕ�R9$g��U=5��_�\HbԄ��Yڳ���>��W�;4 \���uin4���o�H�+ߑ�e��g�ar��H�� Tӽt����9}wd���� ��FG^h` U�" -�G4r)�C�n��)��$T��\�_���Ny���r�����{2!�ϛ]R�	�$�HUq>��k>ɧtn�*@�`�����#��'_����E2n�=�:^H���1��k�g]"YR��0��ͬ\*FT/a�n�z� �����E�������`�"���4+-p,T!��[;�����+����\	��a��n���'��s�X�x�.Xm��?׀>�s�/���ń�]8-bUj��aAd���͟�J#$�A�k<�^zJ�%(7��ϻ��3�*jK0G����HK��������|���6����e�r�(	���K��wHn�]��ƀ�w�.q��r�ҋ��n��H��N��� R�E-�{����;�sU7i-7|�xJi�5֔YH�zH�$!���HS8қ"` �FB���1�����rg[��A��!H�.�Jj�_�_)5�m�7�Gc��*Ƨ�M��!*Xr��*����c�l�9ł>�r�S���Is'ǯ��@�c�P����1�"�2����o���S�w-�H��%��feO~I"��)���;��}� 7��f}S��H"�hV��Pnh����02ڈ}z��G��Q
r�R��m��\���*����������$�J<+�^��~�ng�˵�<��+]��;g�����)<�����	��L�n��X�1r�󫔴��|�T�-�����C����+(͐7�H����Y�'�������O?b���+]p�[�u�s)|� ��2��Άd��G\�Er��v��'�e��ЅU�R�#,r�J�����ڊ�����P�&R�f�EG��7Y�S��1�)�Q��j"!�VK�O���`��3)ʐo���^Sp� �x���$���h*�9�_\�1�\/������l�,�-[#�]�q&9St0g�o7�A�4��0�B�3X�42�^Ur�Mp��*ЫW�e��ε�%����<���	��tr�5-"dj�l�F�zd8�o�z|�v�'E��D�[�]Njs2�(I����匩G���i��-o����)�������$��� ����9u�t<�ahr��V:��2�����߱8;"
q���7��\N�S��í�_�1��ݯy�4L�˃9)�����!Y�2�t��2�tg��`)�?x�+��q�
No��w��|�O���z׈����䤎����s0J _N���'�~2k��~���,eZj'xԂT�Fvo�̛�~�|8�,ca�;�NL�˗I�E��7:��dL���ד{`t;�k����=�d6T?@�w�vg$��DXSTW�yd����;sv��
f��|a^>R�oԹ���!��f����P--B���By�>sҪ�G���l͋���+5�-�n,_oA&�#^��5�x�D�Km*�%�1Ku����w�د�}�l�[^�S;/՛�A�0��;��n��6�0a�0R���@���!Ԙ8�HۮxW{�m���^����b���ư:Y@e���y�N-�"���6f-�:�G�QB������a��}ދ��E������z��51H:�_l�&���9�Rl�B��y�Yl�Oe��è�b�g��1J��f��=e��9	�)�W���Up�.���ȗN�ފ��g��8D_سNs�nω����6��V	Y ]�x��U�&�{~��U���+:�o��<s�)�r�u�.��"���L��Ԍff�i�O����~��(e����?l\��~��A��^��έч���m@Y�r-�v��DH�@�?{��gx�/���>�T^$�P5#��i��n�|`0��g�] ��5#�K��V����nv.q�Ӏ���A���\���E�u�-b������;�k@7�&5��N��w���P;�ĻBU�`�E�@�?粃y�]Ӈ���Y�Ў����2�չ�<V�$/� *;̙��/3$_���u�6q?�	�s�i@��s��ye�g���t�+Q3��/��~ *f�6i����?~�H��qt䄢�ǋ��Ue��A��fS-[mw�?�U��u�O"hj����vx�����
�Ӆz�
!�tj+��(�����T �=!��.k�N�n$;�;�	E����Ց+�1�}6�wt��5Ap&m�%�V�	�B!�@H̳ܢ�ٲQ�!�}8�u+"m/�5F�]��_��ֲ�\�
7p�1�Q�S�c�;p׺��q̈́b���7�Ͳ!����dg;����>��,1{���yI�!�IX�Y,-E\}-hZ��bq'�ٕ�Z[m�s�G&_�r�V!��s�����x%X%S�cA]~+YA8G�`�J�R�V ��- ]�1�����
w��vo�\;�.{�À�k*©��˩yн,��/�9��,_��|e_�96�%hʨ?0�i�)uw(�@h];�([X�u�P�?�H@tp4W6�)����&�ћd]�[�D-^Qv} ����J��|*��QHh�;�0`J�f�R_�	�;���R��Y�r9
�7�39�l*0�tb��;����-l� Į�鹷�"n^X�I�S�4f+��s���}��]�,���~@�Ϣ�teBT�Af;�pC����K���p:Uϑ�^MH�=L����TM+��3�W_��S%�_/��+�=�G��Q{�j���c�R*i#�kv�LG>ۏ�,�H���qÁ��Q������dzCưR<:�hw�� )%�:0g˕j#�0bzFb�<uh�2;��:�c���g��Am�[�)G@F�4����B)1'Zt"��Ac�v��Z���9r6�.�q�Ekf���
��B�����M����.'���$W�������0#�1���r��}?#���<U(�CjsUTuQ3����6w]�{��x�T��ċ��^5�̔��y"ް`����D�v��ƣ �.K��K��	���h?��z�X4�Kx�@�`eYǎkY�o�����R⨂R9�yL�Rv���ޚ��4���$'m:^��f�A�'pR-�lW>��(f���X:8NI^�].�̓M��D*�U1��ߐ-��aUL�u$�I�n7:�G�L�r�=�䰶Ӌw�h �L�F���k�nF�?T��:��.h������
���Gfꌏ_�[� �E�>{��M�g��/?�fįTR��|��G�N��XԀ�@��x�-01�ee>�c�#zsv��f�ӐYDOSz�K6�\���=΅oO�3�!n�1I�;ˈlN��y�/_����VD�'�i��3��<��ũ~�U�h�xU*���No�oG����?�����³(��s.� ����|�4� �,1�RY�����d���5al�(�.+��T�t,�X����n��)���?+�)I'���=xm�y��)�7>�9+m�9ik�:;V���Zt��κ�.�P<BԼ
n��W̽s��>;����
��Ѷ>����ƅ�`G�
̄"�x��럸h-yDֱ�)�����x_9^�"��2�5���8WDr�u�"F+��~�񪢉ث��^6�a�E�׬�ab�8X04���S�9q��r6p�k�����<�rS�n���!�E�A��wb��hz&�S��s�Q��萮����I!�����⧴�I\Ӧ\�� Uy�b`9���q�J�|��x��b�W��~K�7����%�6�b�I�[����޽�:���v�P�O�Z'0&���r�}�A�F�̰68���?�<���x5�Y�=΄�����2s�����7}���k,��]NO��߮Ls�}n�A
?Hs�=_��#�T�.Eа�H�᲼4�!��H_�ڌ��=���O��}��|�KT��e���$bf��<<(Q��%��91����dK�V8d�%�B˗'�?��ʮ�����ݵ d�Vg��I�q�x���~�0t9p�q�+�e��K搇!�}�1�����S�~!����l��%�5�W9W6_�?�C0���Q[t�`s�@ �..`b�z5{	�y�����2d;��N"F�H'�;�8oP����ޛ�`_��L��vu��Af�i�.�	� ��]P/oX�0�'����Ez��P
�RX�K���+Y�˽��a�p��p�җ�{G�U��lz�P0T�^��;e���aX���T�����4Tz�ʪy�45��&���v�?n���[o7�GCJ�8z
��/�=)�=��<mc>) ��q�6�4]�eU.��]/"hغN���)V�� }�s�E>�_�n��Ů����S�c��Q��z.����Xk�13�6�ֱ�J7���c���H�@�_v�ٳO��[�C��6�CE:����*YmϿ�|�ގn�y��[:�Z`��F�о���/��J��rϳ�R.ݱTj�E%�Ash���'H�R]Et҄�z�)!�d8wC����,�?�����;�WM͋+� �Yfڈ���
��)�*�x+i��f�l��?Vǵnk6'�~k�U��O'���I'�R�>�R	���VX��	z,���V�VV
s�u�H�\��%t��L?�
�������Z�a
��=�������-���Q�C.5��p��ܝع���F�Fq+�!�W��A�6�hPj�F
����M2K�٪,�J2P��m!�y�dx��QV�b� ��@��~�j]�ʚ �y���P��d;�f��%�����q��8횠:�N@r*���ܥ��5d�1�d���/�鿩pQ�s��r�t�-��p�_��������H�D�ɐO��A	8�9-�<���#WKpۯ����g���v�0ܮ7�����7B�+f��lRJ����ޖ�{ܤK��
�pGxۡ�ixUv؂�t��V44}�
:�;l�u�������aN�j��n�[��pi�\��V�W0��iI������o��%�ѓؙw���?��#�¹�dx_��^n1�8�aqLas�a�$B��D�\q6oim��+:G\�!�fz��t�B>�����2�LC�G���E�� Ȓ(��*�݌MH��p#a_��T�<�?^M�(�:��#���9�	��Y��-E6rB׆���7CJ���T�=��/�T�C~$���6HH��#	��b�6c�W<��E�S���!j��7�\�g{P{�|��'���{�R�N�h8�#U�n��.���T��|���jp���T�#�o{�^_h�L�f��SV:��r�>��e-�������e�c��}wj�B�Z#�)J��:ʹV��BςQW)����{�|m;��l�(��[áA�Fx�y�݋k��Va��P��;~�7A��!�k�p#z�����1INjc���}�U
,�`�k��R�Y[�U��3���^\�s3G��S�R��D����	 `a3�4P.���?��
�&���D�%����<H#,I�/XPhU0�I!������ǘ3k�qiӆB���-�nw����{u�Ǐ4%G�;*ID$�n�!v�*t-��N�<��i57�b���b��^�ڌ��2���0#X[
A�X���>ϩ��ˇ�'V���j��;���7���w�X��_��p4D`��)~R�F�~$9K���B�� �CjO�>�X�)��u�������3Q��D�u���^��#�!�g����ބ�s�B8E_��SL���)_�P�.s=�&]u���P�c��Ta)�򰲵�fZ�e�Vnͱ����g�3��P��m�c�����a��"X:�E'�@)�4K�����>7�͡���f7��:7��=!���H·轱��^몌���kV��c��P�&�.N�&+3��~uy�ݟ�nX�S7�|ӱ ^�5���G�e�`���t-&RU���<�V��y�k�xI����RuG����`9f�
��ś�7TW)r�7,����~�U�<F�L�rʡ�YG�(e�U"�&S�%�.���d1=�sgG`�IL��o�v�M;��}�@#�O��*�u60���,�S���u�U �ލ�!�&��W����<�?b=c�ޮ:O�()uK�������Z����D��!;�.�'5���B���r	Q�D"�~��ipv��Η�����]�U����]��K��,�m��<�@2����ޕܤ� ��{'�C���	5�@�S����y��t�"s��cNTDvK�Ƀ7AH4��S
�T�Up����;Kx� k�G���j ��2"d���.ʺ����Ø,�h0��)�lT�Υ�@$�D7�A��1io��3-��Q�|f+��V\xg"�ǋ��Z&��un2O�&dU���D��~O�ч�h0�����8;��V�3�������3n��z�EǤ0��N:B�U�\��]K�U0e�-hkc�X�H�CΩ�����m�K�)Ճ�Q�i���ױz���{������ f:��K�oxH�Y��N���!<U�����ws�#47� �G�7i�qG]?	R{A%a^�fe���_˚���;��
�KY�g�H�-�Yj	��K��k��S�?���Ky3XO�|�	���]��d��z��t)�E��-�95�ꪺ��s@o
�y��ZCJx��Ǆ��*?G]�s u�@��ll�)���Ed7N�%T�ݎ]��J�?�F;\�i,i�Q�X���������;�����4U���)^�6c����~w��A|�t�̶ɨ�Ѩl�/GFXi�n�m�$��lp)d���6BP5��\�&N팿ᤏXEgk)W<�pv��ƨﻼ�DQ`��6���N�n�Y����{�k����R��O�\��Q�u���1^"_~6�^f�>������*�{��_{~�U�������m!�6�!\yI����4�c[=e1�Nr��x3Z��/����"��g�WZ�N!��S8���B�4S10�-{}Y�:$��;|VG�>�8�>����gڵ���~ݝ�9ĵFɞ�B�ԋE��F&�5B�w�xb�]h.hx��x|bh�
CM�L�0Ѣ�f���Ck�^�%���=�9?qut�(�]	�e�.<>�=�nf�eS*�2�`�K�fk��Ecu~��J2Ғ���F���ƺp�|��R�\U���[�ypj*��7���Dq.;�^�P`���3op�N�X�b���j����]eoes�ֈ�X�{�BVnx����Ib
�u�2v>
$KQp6�]����螉�ۍ�Q(µhdE���}���2���E�+׬1JK���˲�э�c�6�g{��w[J咳�f�ӯOf%>����x�o%�u43�Cև��_�/���G��65�
��F��,��A�zni0�|��-s^�y���F,�5&d|Wp�����4��jj��X]O����
p�d��-\�6Y?�`�� 7�,����2�nך�ͽ�e����=�AqŁ�����ǐ?X����n��#	��H���?���_���9��A8^���ɲ�*ʚ�~݀W�1���)g�$�m���ܲ���Dǂ	�r��/�1����^����T,g�Mpn�f��I�S�����8��ǥ�Y�dJ<{��ݝ�hIY��w^��E��`H��qM����"qpxg��Yb��"�<�HJ����n�8��.�/���eg�^�(hV�%a��o����b����JYj@stK<�����_@l᱔�?<_��g�����5ݪ%����⁮Z���0�VN Z�f�B�r u5�ݍ�h�42���8
�� z���ϺcLiw_  �!!du��u��nn�< hC�ql�ճ!�����o��p���ܥD��{�y56���9�рs|e��<F. S���S�r�o�_�Yq��l!�����d.�(���d�2�O��)��	�9L��\?e��c�˼<R�$��i~�c���{�D���i3�O��C]�Vs�2Sv��j�߮Î��^Sk�g���޺��O�r����٣f#�c�Z{Cc嘹lmܻ��KT��N+���8E�3 �hv�/P�!����nI��3�_�Y�}=�b0�<� ��Cbr�R�	��6�O�uS�f�4���Ѐ�����5k�k"�Z'�3?��)����Z�z$�<��%�v�.����vq�WQ��X:�ntK�~H �ϻ�>�fB��F%Ք���Srs�y>ۄ���{&�g�����(IyE	�k+W�B�X�^y���H�nUi]JJt��T&�ٖ۫�[�G��#���8 ���ѹ�=� ��m��g�H�zl�Euq��&7y�x��r������� ��ޟ��u�xN�~�9l�c�f�� �Ha��#�|�ŗ�6�w���$�p]<��fy��q�ҭ��%G#��g�^a;��qL��j��:��@d�yn��	tm�e��;���$f˨�s�n���W�2kA�呑�)��A+�mr
fS�!d�N�TŴA�h#��hB{}I��D�|?����6��Ƽ���ԍi-���E�m��qA,��)����	R`��O� �b/_Y���X1�w<Q78�[p����79궒
()�=�݂���i�Җc�`:��'�B9iE�����]�9�i.�^תj��&IӷƢe��ye;�ӕ�K�g���-b"�^��ҁ:2��K�.�6���
'7S�n�}@���%!�2lW�'!0�t.�[�F��\�Զ5������}D��/�Ժ��k`K�w��?{F'���X�t�yg@��"r��|�\r��G�4�"3�`�b�ob�٦c�q��L�3�^vҧ��,��*��Z�u/0��/���E��J%m�Fn
,���{dJ��H�?�q�,
7.��B�K�ݰ
g�N"7��YpBtOM��ȡ��gXe^�4OW� s�iQS�@��
��|��`r����B*K� �<'�&a��y|�՟�D��;	�����\T!�B���T����Z�n��g��G��j�﯄�K��l8�, J�c��-D�W���j��ϋ�
B���Ky�7tF�gil#Va�������i~�S���n��\���@�'���h��K+�$�S�k���5"@83?�L��[�Ж"-8�:���OBےݰҀ!;�$���;���d��ۋ��|�b6NR�W�"`i�<������ZBt�V����
'�ãH�Mo*����F��	q���Z,�&���
a{�_�}!J|L#��q��q!�j�b�@Yy��b�n��pR�]�B �,+���KF��t��Fr��$�S�9�;EŇ��XD��sfp�1�G��%[��]����gm5�6$�}�w�ݖ��?�t�N^�15eA�ź�e��H���Q��c���J�'ss��n���{!�}?4��
�Qp��`Al����=�H �M_K/���x�X�	(r<P�|%�=K�s�s��\���Y�]���́�?Tve~�+Gs�"M����S�kZ`Ej��qAq�,���;�ٿU����8oΪb&Dم��c����Sh��"ycЧ�܆ze�3윚�n�/��5�P�R�vLm�:ͽ3�I�`�B3�^s����6)O��,b)���6}Ywf��2,!<^� /�(鸕�9�Wt�����h�\-r��T��9��[�;�fF(��_w>*�7�X�ɛ��r?&��;?:����l���_*��&Td������U�@��>��g���)=�z���k�Q�S��B,�lc��;�����n{��\�gk�uM��M<�ظ\·�k�\s�￲�=5���R��Z��ɑ`�_��YsNq���+Zh�Q�bڃ7��Gv�2���o�JHc�|9ݏRYӈr���B���>i U�[�S���ՉI�ᶬP����P�Τ�\���ٻm�ҳ��(1�i�?����5����0Ks���X9ח!���,�w�4ՓM7C��⨈��X���U~�Sk����.�Au4]+�4';����j Qj�m��}+i�����r�k���^:w�+et�W�=ӽ�5����`a��%ʌ�����} n�5�Fl��eۂ�l�48A�}�skԤը��-�򍤑)�R���YNB&랖�1��U;
?]��9>AV���_h�Ӟ�G)���B>>�P=+?l���V+�Bur؀1٢���iaEى�e��W���ۻ���̼�y��+x�2�^BD�1��*��P����E=6��x %O/� ��G�ā�3Q?�B�f{;�E�ҥ�Rmj���+Z��BD�8���W�h"Iŉ�cS��W�e�(w2��MI�oi��������h�1�ͭc��02��rߊ�\�֏c��`�U����H=��s���⬤�;b	�POR�hb:���t6'�Ӧ��c�>�Dn��"'�QT��9N��X�-O#8��H:ؿUd���\5q;YG�qF2M���;���܀�i��73�~���{�������� 
���)�������FN�U��^ʗ?�r]^�(ؽ-7�)���;{t9Tq��b�UkDo�D���'w[!��A�kZv�S������z���,%��$����Qj����w�X�O�ٖL����B�����(���%�&@J!-�����ei/9��[H1�\,y�P�D�)��[�o�<s��/�3[�|�����&�i���)hG�4B�#�\ֈ�݂Z
l���*�R�\��|���I�Zq�=���x�Կ���	`�����}�
V�=m���1���W�vH��˶�:������"osk�$� �\�=�����peHبnf���Ì�
Q; 	��~\�u&�N�+M(Bk=X�f=�#%��:0P�����Q��:��P5��Z�9�ű�|�ʸ�������� '�;j}P敿OP2L�ߗ� �g^pb�d����]� ]#c��mr�ж��6��5���o����8O�_��V�mw���Kݠ�u��s�b�X�;S�S2O�9z�(2�$�fԻ4����jۂb�2}r�6��3�=K�~�s=/�,g���,��4Zz������(�fz&�����ͨ>�qk����蕦�o�-�U;�(�;=���$�O�a	��"�.���۽��D�8��ʕ�W��z��E�q�6�~���c�q���#9]�5�R��(�3���Z�%|�5m1'r��+��BM����mD�_-���sV�碏J.�\���#�A��Q��?�O�k��Rr���]nkX}�-`K�$��-\�˘����O��}F�i������x�r6$^8�aHn�-�W7�N��m1z'�_�ֲ�a�]Oe����!�!|�c��GX<�~��������T���F8�(�g�E��#=WQ/b= 9��!]����m'�3
3υ�ڧ�G]`X�_ϒ��m6R�gP�bI{�r(M��z��z��{q���Jx/n�z�Z�~4~T���\����@n��e�a;ͷ�n|PD�\4�2�bu�<>0��t�sp����.�[kF3������F�X TP�4ex��,��+U�� {%/~�����p��$^���Q0�&�Wa�qz�a��(����d�(�޺G]ON��7�̄������V:��d��=iʉ������u����>�O.������[S��5Ӻ����R5͆FN��St>�#[ �s��f$?���<*��}�v(c���G���Ơ���a	/߿�(��H!��FEQ�`��&�"v��{2rG���Ys�+�ݤ� �'������E��`\Td�8�=���8�, f�ERU��["�*���ɽS*����6�����lE����oR��0a��]��+e�z��P�>�k�b��D�����7��in�M1�HtŃ��C'�i^�L6͋��_�˼����3�;<�J�8"�uǧ��5�/W��	�#�.z��X�﫦�~|zWk����}�s�hٴ9u��c����ȟ�K)�B���D�h
����̈��?Y��b0$��+_�Y^���|v�A[Շ�F�����T�.��z0�d*d�_�X@�:�G�n�6I��F[<���^�rx��Ak.� ��n%��Wػ�����m%������U�.;�-^$��F��lͽ��l�?0i#)��Y��/)*FMi!Xe���+�)�������Y�e�"6�wS��w[b�'��@�@�m�C��A��ޟ�o@A�Hd��x�S8�Q�T�g�
�4F�+�.���� ڝ6��D�a}rS ' ��JW��7�.�w�nK<�s�ϭ�y��D�~p�#�D��$�kن��=�qV�����?�W�]����d�3�U��p��^6xa�4���GRX0��� a{59��$���uD�I\s�n�u!�K2�����f�?��d�'�QB���J�Ob�F���`�x��g
��s�}��q�3kպ>孙��E��}?!;8rQ��az�3>HZd��]l���䴏sw�m�SM�G��\ѳ������zE��3�,�ŏ"R��$Dy! j���y��T ��<�����zEVv�C㵣[[���ǇI�7D���w���-�V��P,�K��>��x7����GM)~��\d�c��"F(h�U~�(#KP�Y5#6G�H�T�eK���L�S����>���~˹��8-�����U�jL��]J�� B�f{Ќ�*�!�	p��<ϗ9p�M��b�X1�S�E/�P�$)�v}߁$׸q�\&��.dq��\�OP��_U���l�q�'��~��*���8��?�2�߀A�,4Hy�ڂ�wZԌ��7���W�W�#��5�i~�	
欱[�����G<�!6;2Gg,:A<�d����@d��a��:�m&��ן�E���,�g� �f�,�o���P�Na6�A�l��Gg�Q�I�Dx��/	/`�3wP����y��*��-�/��f����]g��D�<|�5]r��bت 4W��<�~�ZS�������(e-R����������&���q�t#������y�!�3l+W7ʨ�ߘQh>��;��w,!���x������!`�1Q\�<��1Qh��ķ�������7� 58�� gW��zn��~]U�oۄ�R�aS�7�W�[zK���0�!�?��^e�s�/�ė�Q7#̎[�l��y"=��t�=�y!�+��~w]3;�%ǔ��0<j{[p��ɳ-�'-��t��F���
$#b�)���/,h�Y���hVz�,[���D7ܑ�"ݫЭ��H��k-�W�%���Yw���K�{��B\�)
��5M�8�*��/�^�Yx������L�`�����&���K}�[G�_e�qh"|dL|���"�)�?��t��=���4� �ȡ���q�l�}��$W����D�C�HTL�d�lkeEv�zN�z8j�m�P����e�p��Έ�Nz���m��s�~��H��0<Ya���{��G��nBr㠚�#ȍ�S�*��W=qb@vQ�
���g `� M��3t{R���,��O׎�.����% ��j#x"��Y�=z(o��CU��� J��ђ�E�
�+g�'����.Ϗ��RD���n"�yf���9s�ٲ[� ��V�L�0����\Im�v���ab����*�a������J���3Aam"SE��N�Z� ����nb�9KF<��h�޺j2:߁Ģ�.�d�eYݷ�@���J�Zm(��8������6�	�'��BA���#��Y��g������ߛmk�(e�ɿȧ�P�0j9��� �ݶ]���w�S'+Q�)�!�`�vL���m���%x���Nc�9�֖Ŀi�D1E���i��Oa���gD�S��?��xKV3ݶ�}�@���EaZ6�>g<�5p�f;�*N0"�ۖZ��>��<����p.�N��)�׶eee[::�~�o�Ռ�7��[��5�4��Db�ZdO��K�~�=-�!<�^2��A���b��.�
9[)zҡe�i��t1��#�<����u�~�+�������2��kk'A&M`M���M2��1Ghd��k�����<]j^E�.c�V<�q���:�H���m�z�T���cLF���8�������߭9'����m��úXE�\��l53��+ňgf����W�j�K�q�6� 2xRq��5���K*y���g��|��Y!r�Mz����gBJ@
�����>-_K4iIlX�g)��dC��sK�,����d/�!>���l���/����,Wb���`I�%���<E�0=���q�]$�A�-n�lBs�U3��\��c,ޖ$�X/��!N��D]u{LTd����Z�6_ǅu��Ӧ��'�<V�Lq�8��xG������	u�+��<B�xB�V[%��ˋ�S�_��s��֣�*�C%��'�'���%Ǡh������o��Y���\�@#۽|���:5>@��_����r��w�����`w�]�~��>�ך��%l"�(���Ȓqw�k�+�=������'�q�����m1��{�����55(E�-;K��w3Wߔ�����y�C7r��}�'��Z�2?(��	. 7�V�I�ʹ��bL��9�����z~��G�,���b��������p'�hn���AO�ub�D��_����u��*[��;�%5�0(�G�9pc��*||c�ү�7�l��n<�7!!vו\�w3y�w�z��LS�ɷf¬��!`]7<�2cr�-����H�l�ᛁ����T�E,W )���� b�s+̲y�;aR8�3�U}�5<�QU��*���`#>u�]3tG�|�Q[��ݧ�<1]EqxgJz3��nJ ��a�f�ܓ�ߚ�M�͇�e{u���9<��H��{s�P}��R�]ﺹ�|wXp8u��U���<wM�o:@���dgr�	4�{�$Ԕ�ŭFR����g�Ƭ�)�C��&t���t��SU!���.�B�(@�<�Ը���;r_�N��wݿڰ�~J�e�<ru��3�G��P
&�����p ��r���N�/i��1���<�^Cl�E�`�LE�)�R:�.���p!2��Ε	��Ռ~v�"�N��<FvEz5���2p�����u�쾟Ks@�D-�Զ�c.��)0���p>���ψ�'_� �r�-K�)ᅩ���'��U����vN�� Ɨvo���;���i�ܰ~��$��Q�d����@f?��,�S"S#�Õf���v�=�g:��v��q9}1�|��,�;�ӓ�#�bDe8-g�_v32�c��ݢ�P��j|5���ū<���V��)Fo`�I&*�_�6�}�P�_-�	p����}�D�־&�6S�{P
�Y����b#���Ȳ�,tx�Ɋ<i�Z�,�i�����*ޓ]�^�{ס�ɿ���./�jydv�1bu2$vֶ���"�q=�,�6���Η�H�X'�S���t;ٓ���:���^�r7�wTJ쉎&I��}>�>rF���~c��$�yj�,��h˕5s��ƚC���:)\%���2^�i�p�b����1���Hܧ�e�y��$.����7z,����Dtc"��G�ܫҔ�ܽ�a.=��h�����Q���Ǹ�θ�ӎ���Q��t{n���k�L� ��E������)
>SM��^���F�l�J5<iF�<���H��.O#ᵕ�ms�*�W�V2���u��Q�P��4x	���p��:�kvϼR�)W��t%�/�)�'����k�p�栓���a�f"!֤im�~�KB0�E�|��EQWHQ\S"|}�n���� �ρ�?�ʽRطU�1疠�\���;������_�c��A
Ge�`p/`�g��䍍�)Jq�vl, �myP��@���� ��
��<��(P�Qww�$j�����/ђ$��o��8����
���V�)xB����[}Q_pب���ҳ`�6/�,�Ѣ�X #����!w�*���"R;K_�� w�afmyp#���Yr��Egjj�������*չ�ø
��`�?<�������H	��ḛ@�Za��`��iyW�:7=9�cg_2V��t&3F��E�:�_Q�M X��{�#�KBU���;�ܣ��:��ťI%}C�j�~��'G���T�g�Y��<�x�I�����Ճt|������g�9�_���䕨G?��ŉ�o�j���7����z
��.�wPLe�9��泺�l���E�n0)�𫀒j�δ�'a?rˍ��HIn�C��~�F�������I��n���Xe"�s*���_q_��`"��UJj`��{�[1�7J<l%�U��p4�i����s�a�B�E�n;��u~��׈а�\��Y&��C�S׺�=W���2P�Ҕ3^c���/;ɨ%�X�h�v��N.*��6&-v�jo���v�_�_�]��>����9_��u�2�V:�6��~-���A�/����O��A@�LQ����y���Z���:��@]��E����D��F���4����|���d�r[�%���B6m���ުt�D�韠%6���n��`,��i^���s'V���y�� AFH��,���=�4��R�k�<�y��\H�t�����ȱ��|̕Q�BFF��}��ߜ_�~���\`�֟S0[�Cxz{|r�k�I#�LM56��z"[����o�7��A��0Jb��ɷ=�-Msso;��^f�	�V�ec�s H�>��K�QoR)���%+2E����jE	>w[������n?�v/O��l���K8��s���똃bf���E@-��h>|T��
^��9����!Z��|��j�Q5<�P̈P���KԀ:�`C�d^q��2�Y�΁߁j+I�(LuR������E�A��;�-J���|;��0�ƞ`w��%�$ �͸�Vc����X���p:	�G���^�kS[��jSd�.��f̴fWrʷ��),���!`KC˛��F}��� @I��&����G�ʒ��*�q���� $�!��5h��'Mn{�פM��*���T���,���/nfI��~������������c����)������h.{�j�շ�4�A�q0�nN�-o\A�mp�L�#��Lx�
&�ƃX��KUI/~q\A��1[�@x^���z���=���+��:�V񆃸2��<�ӷ��]t�xpW;�|~�<�����^����=��@Z�'�2Ű_�����w�ܶW ����x����_@��7x�)4R�h�k�=�b!����9.u����ďn�w���k&p�[2_�IRZq7��K��w)d��B�5<ʸ����aCcG�!W>\<���<�?���_��
{ۤz2���h�����m@�����b.��eZ���A��P�^^�g�3]M6��B%�-��K���.4p�zvS��}�nM�3}U�N���r�$�a�58sN;�
EE�S�7�0�a'�p|���(��!h�ު��l;zy牏�%�X��K�r�3�^�!��R��d���/�	�Ńv��K���!��T�r_���p���%�N�>c=�I(�HJɩn�$_���;H����\��Uڭ�x_NiK��m硞%,\�Gʊ�H�� �F���w���iq�Y<��P��V`�����l����a]I�q���W4����������)���њ䋄]�pF����	Cg?�KCT2C瘀x(Ż��.1l�yL�E"�@�����v Nj5,tI��*��F4�a�p��-�=�5o��9�&7�պҪ{ޔcbH��z��9('�X��6ȫ|���l>te3<jeDWG:��v��WS��b
?Z&U<�b�73�2ЎX@���������d�i=)\�Q��l�Q�*:�=~	����U�bǷO�;�${�WJOR� '��.Z�r�6}��W��i%�n{ҟ����v��%m�T�r�m#%��_�`>ֿ��e��I��,��R�y\	>���#oP0?�ׅ�Πk>�����H@�t,=�����n!�~~�d����H3"9?mqU �eM��2��6���0��<Dr�]Ȯk�0�m�+���H(�Qdb���E������!@;*�m�L��4%�
]��!準��G[:�#��d���"1�_u�����6۱o،�.�Y�Kر��L�F��:�Y��E���E̫�I�k��ks+��+٢&�¨��Ph�[-8	�5������ȏ�+��~����.{R{r�N�e��TĦ}�آ��Y���ыٷ�r�"�|�|�t��=��s8��T��y�f`��ب�M��Y0j����>��AR�`��w����N���S�#���2q]5�
i��Xf\�	DU\�-g��'�.����C-T/|�,�^��U�q��Yc�p-&i�-Z�Tؑ|]�h��uN�!l�u^�!ݍ����$c����wuI������+°�o��P���|�-�������hZ+���H�r����>�*���:���I��(�(]�c��_	1�h���ڶN�j���*�b�5E�����K�AD�g��s��rS<j�&����ku^����zWr���fg��Yi�s	��k',�-��,��ҟ�݋	��nD�Z!�@=�5a����,b�9��S�rƖ�t#� �Qs�1hI���s2��O��fմ�+� �1��7��/�}���mt�}݀o�
k0{�Wn�ox�[�q���AR��IJ�_�����8{����R�-��,Ы�8ၣ�[̿�Zhу����E�ki�������U�4�,���=#_�n@nb�n�� W�I��B��d����J���\i�_ϑ�A�׼�
\������f�\��ť%�ƽ�-���Y�:���ot��Ȋ��m �+\��~�"�OpY�N�y�f���h�v�?;ބT<
�9T��b;M5����Ƈ�kY}'H��[�xR<��[��T1�~�����Rץ�zh����I�V�2��p#�x� ��Y˥TJ�|�bb�Zf�#P����l�cSu��Õ�<���F�nAN#uo�Sx�H��H��������K+�186����vʨ8��3���eDkj��F�c-�.�
|h�ELu��ɖ 3�DLtY�X%s^Ȁ,��,/�f�TYTWR'^��ky=���yK	S��� pv�'����]h�T�k:.gq��D�B����C��UϞ /�ud����i&����i�w�����p�G��,�@��-�gސ ��I�!B�yr�=]Ik�g�X��\���\1\�����c�u�v*�f �ҰI%��2�V��3 l9SĿ}*�1fe���r���7Dh�r�=�&�9b)��]��<��f���%��`�+x�R�V��c/�X�@�7���^̜⼩y��F��6��L�7��=�[)E	���{���"x��
�ZG�;���~S	g����#c����|�r�0�f��>J��������5�����\�g�K�?m�(���y�/��匝^�>�ݾ�+&� ��na"�+2:���g�̗feO�jͦEDO|A8@I�ȸR�e�M41(K���|�o'��T�vC��=�ʕ9���i*/���������ce�EB�Ո B]�(�#�޶&��p����~��;-�tD�+I�t�Mp�q�m��c�j��0>V�h�&�����K}g�7a��i>��>D�O=�Fr���+JفbEQ�`�9��o��w����6��5��|��,��"[p6Q_��$��n`�jVUc!R_��/K�s��pI�S�9l,�'@F�P�����,��b]�'��ɾ1�c�ag�ŀ��^�V��|�2[������B�}U���,N,�cwDCLښ5�2�0G �9M�A_MƩ��'��B���]{������_)��򩮞�ݬ�y�(3�=�	@���=E��π����_�Z/=�C� ��r,�/������A�ITQ
�C���:O�d���c�날�4�{ 7P�F���+�\v'p���}��p�M���bQ�-�{���AC�t���T�>��b���yau��u�ȷ?l���d����p��U#�����Y�5�x��2�S�|�|���*yi�B3��A��kK��׮Z���T�0^�H�
U�A�O���;�yJj+ո�'a'W
��b
�A;�:��p���
� ����s��0�9��Q�]�~�5�pgԖ�d��f�W��e�hb��>�Ec�I�TooN~���8�]0-�7�:i`ǎ��uEL��#l-,����T�Y�$����3���rR@*�	���o9Y<�1�pM�P�^y~d�P\�]�whZg��8���Ȱz-���u�U�QEW���ﳃAi�^�_�=�8sJ7IK{��S�H9�oo���e�W( �:�zJ|�1�|��Z�J��a�߲�T�T�߅ �+]�ӯ�I]���L8݁�_9Z����2�v2�kYN���X'W5��,o��u�x|�y s�`�eDf��R���z!�n�W�}��[	N�b_W�E�zȴ�H��(�z�۪�#!�"�05f��m[��&����f�p#�����Sz��������)���hT���q�#\!(��24�b�p�@���C|2�+|˔Jc��Z����U;F4=�5i3�L[A�ߤ�P	6�CaV���F�g�I���v&�q�D�$���/�́�F9r��m]G��q\G]�5��,�X5����N({�U��O���XgN��L�2�\�t9�P2[��9yP2^�M�v��b��i�L��2`�3����ϭ��Y-�ӣ[%�����r}=��e��zw�9U��B�>�3�^e��������b�6z�;��ӽ  >@��z�5�=s�Y�F?���^���ز�0�:�Y~�"_4ϋ�f����w�0�8�+����=g�?���"dR[���m�fH��㈛��3Y�ܙ��8�Tnl�q#�S*�-�~g{���Kŀ���= �+>PٜT�����*"�,���r)e�)G��\;�饍h������y����3}�>���7���"܌^y@m��~h$�A��Po�0������0��)��MsG��A�_�<"%����������9`���?�$�CΔ�v�k�&n�u�i�����}x�*/Y0���+�����y�s�*԰��4���)��q���oh�
�n���0�?<I�u�����[� �x�!�V��U��Pm�G���:|���ĢS�u=���u�@�����[偞󖠾O��}=JR:<*�)�C��>�"�"��ׄl���C�N���f)%��T��د����U� �cK$yK�3��𛊣6���;e�6p�W��J[�W��;�k1���^5m�П�Ӿ4�$�I��х�O�] 5*4�_��-]&�~�ʻ\�nx!�oP.��d����K�di��{o����5�%��B�gA���M���w�@����\M��[Mw�x��gG�}��iV�NVv��ҵ�Za����it��m�A��V�c�oG��m���+��[�4J,8{Gd<b�3|֒@t��nbpV���l,=������}Y�jp�j쪙����fX�E#�G���=dF2��E���Aa�0De�f0�p����ʞ!�R�W��S �հ�b#���+?����1Ē���013J���,a�I(T#�����͖o
�[!	��N�8�g���qk\�Bl�ԚL��}0�Ue�Vг�6Z�@}R��΅���9�1Leo���<�_��苼t8G�\`��z�ܔӘ��vp�֓��p�-��|��
�O<�$"8sJ��5BM�V�����������G����=	��'���\�$�įyL_D/�Q�X�i%��u+��X�#�W�8#����c�%���ߐ�>>�Kg\p��l���ѷ�~��s]6S&��������0)����
��9�OB��y�s�~G�o�'���(���9�(D���R�x�r415ק�Rɺ����
�ᓜA� �?QgBOX��e��J��V�y�2M�;%���
�ԉRS�2`��V/q�������9f��ޞ�:�B=��,G8��&�����/I_0[�����Кw��N�q㽓H�Wt������n�5�8�N*/G��v/8ֈ1L�>�����[��cYu5��,���|6�u�%t�\��/�U��"z(�+:$���w��<I@/����/)�p5!B�͈���\�:�L�>P��-Զk�yŰx��*':�$_�shO�o�������j�;A5!J&Dc�e'�%FϓLh���f�p�A|��/�_]ĥ�yI��¬50/d�
��f+��O�&��:��2[YJƏj�����Ѻ/$(�G��v��*�M���������s'D����^o٣Ì:�q@�K��Y�f?�IL�]����v��_o�j�V��K9.0��{x���:���}FW0N_$Gm9�������̰�ĭ�` /)�i!��
�b�#3:xqz���@P��"��b�%d'I��d�'d	����@��B������@
�P��Xkw�)�m���h>�4��Y��N:�&׊���G��/iP���g���y�}m[1��u��W�B�(LӍU`��RQ��ڶg>-�CXӛ/�{�?��͠�0f�����N��rc�����~���!��1�8��9ע�I��+�J�J��Hf�}x�
�u�L�y�5'O�~��u��L|k5\T�RΛ���T����,5�̦�{�w��F�5��'"��BA��u���n� K�� ��2Q����P��#1�U�߮$�1�>v���x�!��f7h�L]0BL+�t�a4��ގ�_#�=�Nz��q���C�5vu�0����}v|�s���~�{c�>�����Z�j$��1��(WFv��[���	�-���}wS�$�N� �8j#�9�����ӹ3�B�;ݡ<�N�/��$������a�U8�B}�y�����e�z��[j@�dyøI�v���N����,<8��1����h�l�X\�R��q?���A�/K��Cp0k,��y�w��lG�5'� 키�I0'�_6K���M� Xe˵�T{�B��tԜ�Ёu������[���F��1zĩ��RZq*���!��O>��Nɾ��7C HZ�q���t���U�E��+��0�'$�&O���Pr,�r}�t+Y��,$�L�r~��,sl��<���tu��:/6��w�F=^	;XK2��$�Ӑ��B�3�9�Kg��0Jn�EX�R�=_�ټGs��&h�.g �_�}}�\ƶ#+��u�;��\����~ZLh��#z��g���|��J�7Q��mE���gI{rRe@�
~��Q��c���đ6��'�x�gTl�SE!�c��4V\JU�5G�A���!�3e�#!�P{p�Fϔ����	�8lCh&&|�-B�:�_� �z}���v\Д
q R������=X0{��99.B9��-�#�q�_���Wоw��u�Ԡ#��t	�ˊ�*���]AoB�#�wJ?)$Ԯ��^XC��t�?�u_uB�vk�� ޿g�Kx�	�{�R�;:5-G$����ɔe�AN9M��`�U�N��%�A@�r��I�ގ���� �}�
.�3�s���ێ��H�x��e�M�2˨{|Y����2��s����ɷ+�~6<���.�U0��q�WQ+Y�z9C���^��[���$�_����V�E����OM�ӎ��+Vx͓��H����xĀ�06�2�;	R�[���S����M��ݣ�����,���w���c����m��Dmݝ��a8�G>fĭ� ��Bl_F�5t��b_�T�?}Qy�~����9@��I���C���V���N���r���H�=�u�(��G����!��6�did�R�[2�����_h/*7<`(�Ξi5&�t�g�_+�2�}M�I7�`����w��P	��{L����9���̃W8�a�_�-�������e�(�V�آ��Ev'�8#��U�OFPIN�tm��H/�udy���o�X�i?|���y׾@l��aOm|i�V+��7%n���/9=A�;�K�mm��qy+���Z��	g#�s��eE �=P9\�7KChKN�.���.~Z�ȑ�ƛ=	+.Y�+���D4����u0�p� B#�T�n��ኽF�s�v5«���������\�#�1���>�	=.k�8^�����0H��؛[̍� 3��T:��*�j��+{�C����=��!=�z��^7/�	��b���l�<4鲘�{�3��R�;��i����5��F�O	��q���ʒ��v6.1�P�g�O�h8���'�]�^w&�g��ީ�&�ђ���?Pvyfc��!w�C�j&o�%��,�0�)|��;�р����r���؄Yt+�f`�D��w~V���Yj��N���|2=}o�d�5���H�ߕ}={t�=9P Ih�{������LA���Pf�����1������Rt����&��Pw�+����*�P}��$j~�o�T�Kv�t�WP�	+���#M/��rs�
�?i��K0&ǝ��{��fձZ/t�ǲ�:�l�<Ĩc�X�R!�"}��������m'5yO��;�¤T������2\�~�:�!G���,�Ll��v챇 �	�L]B�ኩ��ar�#� �(F@�p�߸B#�����g)����Y��a��zBGx�f��c��g��<]�pzm�G��S�R�f:�ˁ
����L�&7K$�[>*-:3�?���'������1�d� (�ꕜ�6Z\��/�j|")e�a����Y��S.:�T���'��R����֔���=�nlmM�w��S6�d��0u��`��%�B�;��mz�!�aC�2y�C�m����:phh��|���e����Q�N6��,0 ^�M`S��O�k�ܜ���
ujӐC#/Gkp~f�?��Sp�׻M�ҁ��V�ܐ��73՚�zWp��W����$[q�1�_��(�@�B"�wUdl�7D�M�6�a���'@�[	�W34��0�����W��򮹰BE���AÔy�oJA;�`K�{ۦCd�ܓ���Y|��~Pp�.����*��|����,�ON�!�|(FqP&2������rb�|n�.|f �mJUG�x(��x	CdT�(X<ޕ��NmTR*��S�#R���6�/ĭǪ�w��%��Q���=�d~�B�*cv�0k���t��0jѼތ(��1�{�K'��	�}��r5i��S�v��ڕ���D�$��#PQ�w2d.a�'����ڠ��^�^��f����TX��\�s맑Kf�{�bF|Ux���c��Y!˦��W�#��ո9��p�M�*�t��Θ&�U=���|V�!a�����֠�#����]2�S)Zx~�a1�\�p���7�����~^��S86c���h�'|S�-�Etɻr�z��a�wA-tc�N �^܊�9�4�]�)�]j�����r���	Ʋ���_�� l���2ui2@bk	��e��C�(����ᫌx����
H����qZƿ�V૔��j*!���t@�k�>�{T4����6�~o�
?�2sIw��;��0��5�Y�ޠ�~y=��d9A ; �T����1�/N�Ò8��(T:���V���:*�͗��������,}���jĵc��ԩw$�O�����7�L��6vc&ԙb�%"q��Ӄ��z�^O��m {�h:�:��펳��E�iV{�Qu�	x���_I���vXÜ�8Z�ת��~f�"bč�v����U�1�Q	�(e��a�)��
�!��[c`5���c@"[`?��!C>��\8d3��+�Q�j˟��
�']Yq�.`�ݲW��,����~����`m�L>F����DE4�����R÷M�kk��{4����D�/��\�;�h]��r�{��w�5����˼6����t+8��*�N���TI��K�bZ���2*�����E���@-滷�Hf�L;��
�p�����j5������|�B�m߶=���F��Rc�2��Mm�u� ���{�պ�k鏡��Kt�P3hu���T��#}u ��r]$.����k�Gy��(������'����-�-�v��'G���+[%�I*��3�zv�H�5s���k�A-�M!��S�6�W�=�C��:g���arO}�3�|{ܢZ{���/2Ud�0�=�Z�΢,���!tCH�� �~��.�)K`<-�]y�K�Eu��޻�+Yv�y1�Y�����)��� �Y�2"6�2����\��b����P�n�����c
+���ZjL�Q���Ӡ���������c�w�&�>�p�g�Z��|��b�	Ӎ�e�QA�v��\���B,��]m��h��(L��_����`/�M�Fڛ��������\M�c.D�(R����@� ���sq;�b^T?�>�%��O.M*:^	�L�r&�n:"���TX�;��� �w��v�8�A���W�9�(��<
��������,�fl{�_�f��8#0��q���a��ܿU�!�jFݍ����
�Nua�Z�qK� ��?�_�6w��v�FЇ��X�Ѕ7:l�k����ȋ����ٔ�-�����{�*� e4�F�1;0N�q���q��$d��#&IGt�*�1����C��ڔdQ-�iJ��Kz�
_���珦�F��J�UY��׭�.S��E�����A�q ��j�Y@��	�����T�/���Ӟ�E�r�Xu��}4�\��M6Ɇ�a��uш ��&�t�y�áչ,�����hH
]w��oM^}�����!�%���Ui	!�Mr(H�e l���7�>���}�����-Nr�C��,#�w���Eo��K��y���h�<��B�;d4J�	�#��4]D���ˮa�=�j�?_\�.�i��z^�\%�D����/���.������j:_��d�"�	�_�:�P�*��@��'*�sɮ̵WiѪa�ii�~�ܒaݒza�/�Yy�A=@���O���&?!����%�oX��랚r����5e�)�w|�x������J�S����W Os��L��V�(_Ւ�v;�t$�Pjv ao�B��@��(�@z�Ϊ8WY֟s]�� pl�~�	_6O]KGf}ȗ>͔Z5��4�^�ib��K�N/zZA����1��D��3�Z���XQh?��L���|�^�{�d4���5���Ȭ��Ƞ��J,�t�(�fM"��|�S|-e�.����IOU6D�Gv�0f:2T����GF?������!��>�O�k��R��๴�>Z�H5�|[TK��?�i���q�ISnE���5or�q	�ѱ����j�=P Nd�� nʴ
˭?5�1^$ ���ݠ��1��cF�
�o@��L�qK,7���ZN5�Lȡ��;n��0:i1�q�u7��$5��lq�e������ne>I�
p$>Xnvw��5� �.��[�*V����4Rd0��6b���zay�IK�.�93SH�'k"����Q��Z�����~�j�T!���������윺C��=� G����毲0��r��r��/G�	|�	��]q�{)�ߞ�-�m+��!�)�wd��h"I|�Ё��ܴ��Sq$�+%���\�Ԯ'J?�q$o�O�V-`�>S48v�p�s����i�`��9i���A-��9�4�{x�%�:��L����}�T��H�!k�G`�~����ڑ� �)�]+��9y�4&�f)	!����L�f_�=�6��*����C�i�\e��� nj���ۓ��3K%�Z���������8V���p�yI��G�$U7���������*i��ל�D��1A�o�Z��\`x'
�ch��@�&"���j��VU�0�@w`��5n����QQ���L����>�b&���[�Q�+0���3�DQ�O�ٚ5\6`��ȭV�֞�K��e�3�U"���Y��V
�o��Ʋ�2'�`�9���&"uZK<T�yG��w�w(���fx|���,f`���?���Sc�*��-�&�VP�Qe%u=S����L�<X��$2�$�"�
�c~�`���4h���A�/�l�M���d��t�Ц�x$�G�i�%���"��V���s|p�����K��2��*t(da�^kv����=���:��}7[Qh�H�楸��Q#�~��c�J�o�?॒������#'-�[�y�ZA�C�!�_|�'F��~iH��seܔ��j](J�R�D*�D
��^kQ�^8bX�φ�|�TO�!>%��aUc��A�ۄ)�l/���#�$E�&.�K(_m	3���dc�9E>=�D	��z�3��_!M[Q���^c6d���� �GI:XĩK���"�z�C�.�뼫�M:t��!�����µc�3�U$�����Oa���N�Q@<�7�����wI.�K����ܦ�.���?�Rl�'}!U�{-���T���i�	�6��h������= 1�چ�q�S�5��D��倮����د�dx%I}`)u)�߿"�M7��u�$��f��+j�nK$�id]s*y0;��po��T�U'�1K��d�)�=;lpR�bݒ����5Xc����t�,�2~фu�L����9�Q\#����(A�y[кkZ[aWo�	��Y�%����Y/y
[3�p��qi}�o����/�UT<���g#�ZZ=��Í�8(D��FCð1��u"���u��N-�y��6D
����F	��K�$��8��p����[v�k��I:P��h�55�L�b��N#8Y�
�4E,A�m����D:Lm�<v��pn��2�5
��
\ٔ�X�͵��1ps�d�0�gţN�Boˬ�L5@)P)])φ�|��Ɗ�(v]�xP���^�u~�:�U�[�̀3A��<����ַ�E�i�ʤ#�IJ��7*�Yx3W!����lKͦ.�űz4�͑�D��3��D��.}xMD���Z'���|&��1bR��7�D�6���͕'��x[���V����@��M(�'���I���l����zC���H�8-C+�A����� �W��Rj����n=�шm�fq�SVo�0�k.�6o��Se�H�]��:���'���eֻ��	����W��@4!�fS{}t�I�:��4j�%�(��<�
Whc:�&��ɦ����Q`|������$�/n�;3]_��"�͋=E�yt��3\�9fOe�\�TA
e\�{W3���ܘY�]�Z�`Yrx����,Ԙ�1�ܖ��S𜿁P�~1�$<���9�	LA�Iu3ͫ�~��o�+-[�������a)j�شI>�bB�G',;�ڃ]yPj������n�\J��D�?�"���z1N��&kk�>�l�L�l�|��m.��1!�0
�3�0`�OȪ��e�?��]\ڍ���g�Q�6x^��G�0ł���~��O$���V�'�(�B_۠�� ��Y:�����G^2<�����oE��e�_�9G��##x��3�Kб��RF�%�i���h��M��8����`Ш��/l�N�ؤ6�����luO+�
�t�ۡ'(���ĥAդ{�U\�{��ص�M�QE�'��R3��� `b'�T�ߩ&��� ��B>�6�������m���%e	�A�h�%�'���hC�m�|��b�?#���=���B��v��!�v9*�n�ӎ�p�$m'��۴ip����%�"�.o�����72ڰB�L)�I�@w>�K�c�ryN�nf��駑y����Nwn������\!��	��Vl]��A�l�"��RQd:�{৤{�#��5�.�����jY����}AWRiSj���,�J�z�Ʌ���y8ai0(�X���!�9}��EPV3=�t~G]y�\��C�����|z�x�Go7ݡ7�ai3i��X��;�^�����`)�H�z}b/H���" �.�]�AY�b]�v�d�S��1���m���}7�,�Vï2j��[��9b)�6*�o�"DD����BYZ�׬���U�f3��`���	4��8���f;�2[w�8����_�*�^��Q�Èo4b>��S�-o�8�5?,���`,�.>������3���Ug����T�g�Ŵ8���2C��(��[��B �7]�voєղ@��q��	����������(�663�%�[g���w�?3�A4�nJ���xLt�N&ˍ�Lp��I�����].S��6�)[^��F~&�:z�+.�
觙�v��w�2E͸P2ҽ���Z\*�rM�T �����&UA<�����$�s�g*J�.U��m�"�t>����IՕ�r���7����a�齺h���_�Q�F�i�\:J��{QU}a�,�l�s'�����@����BD C0�M��Z<��[I��K�K����8f��y˓`�WH�!�X ��hCb/MQ�	�\&��m�Hrà&3��E�L�avT쓡J=)����G��!jʙX�����1���ҏ�U�L)5|�P����Q��˅��߶�:v�5:��~�I;I��w�u�ڢ��y��3	~H���g��ݕ5��(��֥�H�z��88{�d�y
�NG�u|h�0�K�b�% mRGPe�#c&��+���^�հm|��o�6�<��i���"e�XSAq�%��R��-�i0����٠��x& LA�ϵ!�b/a�eU�)\F;"�q�8��A�Z&.�/�c�wힺI)��v��zj���&p'���Y����+�4�	k�-t=�H��P�eFsTM��m��J����=��c���Ȝ��s�l��6`Q�����'2z����PӘ�o'P{KH�:J�>��*�� ��K`N�,՞�����6�	�og}�^�q�?:�����ff�kf�ܝ��<�e�4WP�f��d}2Q�j�rc�o)V�b��3�����)�W_a����׊�-X:�m`3k��CnI�U&���i!6����?ܲjCТ�_�Y��]�ǠP�&�ɇ���tc���J��X�ԥ�����qZ�6��l]ޝ�[�ı����T�vG��냷qќ%$���#w:<u�yN�4�l���J_|�.��NP<nw$?�^��vVF�Ϊ����L���C��}Ϩ^�������=�cN�³�LTj��	�2��#�Ϩt���aZ*2��k��W��-����@(v�t�Y����g�I���ūnǺ�a�=Z+��bX��{ b켔���.��;0�,�W��a yIR��8���|+�d����h�2�2`L���4ᆗ���4o��ƣ���-�k���&�?~�+�?+��'Ro�Fgpz0��V�94�~S�� 6ZM/��F�]^��[Z����Z`���n�j0�#9l�7��JL���6j�<��ݤ�eU�xڞ�Q0��������];�A�+aq����'��[S��r��A�b���'OU�]�"+�s[�ǅ������ �7Ġ6R,���TaʦDІ�����qSs��D��U�ğ[z�h:I)��z1�9������b�"=�h�ҽ֤�*w8�|�G����u�9�~����SW���/�@��3-�Z���U�;���@.~ʤW?~� t�c��Az�[��ڞv��[��l�<�zx�X�vAD��LyC=4����?6�H9HE�T���s��9�pn�o~TH����D�,�eq%��S�G/�K܆��-�_d�9H̛����~�X��WdB�����`Z�=Jٕ��PqʲC�@ �^��\$ys�+�Jt�Tһ�%k��Y,R9~=�[�j��w6O�	<R5��H�}���E��㯗����~�m�7�����S@
�{'6��_D��\�k��p�;R
uzG5�/P����#HmQ���o-���](h�bcr���f��
d��U�lk���$�������K.����٭r�]N��ϥ*��͙��X`�䴐��J,�|���^߽�σF�3B���:�d��D2�ɕa�����LO���h/&nt�T����m�AS�Xg^�:�����'?�����,E�����s/�h��X��,�L���:+	�⎋�k�{z�Zg#�%0G�>*��V���;�`z��B�q�c��m~O�4|�w�-}L:��]�
�nMr�[��E	�s �g�O���[��{(��ϯ�&���u��'��K��]�i�PEt�hT��C�io����+4�h螸��'\��4DP� f!���D��M�.�ݧ���ˆ���y&ӡ6��Q�{H���e5��L�]%�8;�Om��[��)֎�ئ=�+M�B�fI����"kݏs�g~vj���*!�ɧN�����st?��h�����5ݫ���YZ�0�-	�J�X)������7.M$�Z8�`����?	��8q��ƒzD~i�����d@m��	z�#G1�`�SOy�PQ[*u����eտ�z����)��dN��[�l�E��yv�^�s#�NGR�ц~L����qO�4����ᙾ�\���e
�ӬT�L�_�����@��c���cǄ��K�]����?�N�7t-�ʪ���-ދ���	�	�Ȓ���XIfN���H�dP�h\�kӮ��c'��ȼ�3]����h�;���y�dQ���V%%TϬ�܏�Z�������)��F#�yI;���'�2�[�y\��;��&Y�f��#4�p��{�AH��?��CH��`@ѡ3�ف��Q�KvF�A��EW���N=�_�af�>
��n�� �S����+��/�b)/���o+9�|d}�smر@�*�\����}|�U%�����q��uw���{��!���9yF��u`�1g#+(}X�IR���=��~����z����O�lp<�u74X
��)q9aQ�����_���)�����r{�:l�k�B�=�2�΃���"��Β=q��L`h��6��j}�$B��v:����*pr$�6��=��.���Q�|`�~��`Q�r��]��gCKmڭl�Ζj��O�e��������u�J����Qx��4��u��+��(O]��	��_;ln!�����s�y�׿]$��S��q/�ri�_=�e%e��d%�����ބQ��y�٫�d%x�﹧�����춗��=;�)����2|!)�?����,�3܋�Ȅ����ej#٫����	 �^�.�.�hM8�R����?�{�+��p�ϺJz�=隼�Y��1��<�~X�G���s�� �s� 8�H7��||{��MN�,��%�4P�Ғx������9+�'���
%����#<L��>77�ĞJ����WY%L��5���J��2s��`֐+�o���BQ�}"�KA%�	��G���p �pv��!9�Ǥu?W7)��V��[���!�1�z܌Yjݬm���Χ�m��NV�r�eO���1��iw��l�1�\%���.�SNs���jp�2E��W��P��b��_�z��9[GZ+�*O~7#s"��sp���>�v���i	t?�h��нq�+V&ʲ��4ciEN�?s��iŰ ����#��-�ږ����<��9Ej�݊����t������f	RS���U�\L���$<��6�O��]��lJj	b��w�����C��,qw�={cm��E�gi����/�n�K�`Zp #�B�.CZԤH]F�����T؞1��Y��[m��6�,R(v�nu4c��wm�;f3�,��<��|2����ɐM��gv \t���sH�;]B���&�u��a{�-wʏ�_-�(���R�Hꀍu�&,�����6�'Ǽ�7�ϯ5�/����ltj�)#65�D�������`V��K�C�sِP5����;����(�-h�r�	��dd�gl�	1����R���_©`������(|��P���?�W�5�|>�%��
�o�.K�����I��4���3��������&� ����iY1}=�*�V��/Y�ȷ��9dw�����Τ7�zp����B�߸�M+r���E[�����젧�,F4�Cd?�$%Q�.,��V��V��Ȝ�����o�:բ�-'�x��|��/�q����r��6w=�*1��";+ib��ɛ�t�}G��K�a�&E����35|��hs#����z���O�:o#l�'j>�[+� u�	x
��MƬ?�p��a�O�c����d���h�3�}ߎi���)���5��"@qQ�yb���t�'��Ef����F�]b)�E_d�ߖ�Ll�T�}W� tu���Á�c�74�I�t�X�؁��s�C83�:=�I��;ā_iL$��v�_uo$j;v��̱�������7�q�+�-z�a�[<�R���! ����ʈV��]���OP�B~�2l���Uf�魣��AN0'����
�D��c+��*u�B
RN0ډ� �'Dqz;�
*���Y��5*��u)��ﰉ�=���.-����!��򋙼���	К?�������(T���d��[�GCb�VM|'
��S-�Db�4�~�=�{���K��nbɥ�~PLgW�]��W�����p��|8U=�C����EMoyj:;��e���-sH_M_��O�><xb��蒳%��j�E��&����=�XXعy�֠4�
|΍��"�c�� )�1�Bv)4�p�x���׀��?�Q�ቨ�`@�x2�c6��<��_�T�ML�lO�#:�܏�[��I�(�-���gJ�ږ���ㇵZn�H9�,���=-�t��C:���)]P�Q�D�c��`�WP��d�:ҙ����*Ê�P�k�4��e���~i*��,g����\����7��?{(v�\���׳ը_x]g�e�?�>��Ε��Bjk�m��ݏ�� m*!;�v�趙�+��fD���U��{F�b=�K��u��$֯`��5�g��R�A�w��=ccC�5g�9�
�����o�醇|���3S�&�C�ǣ���m����z4�⻴t��R��
��-59l�~�O�ީ4@���//<<�V$���
��Aͻ�
��64:�B'u(�/KQ1?�	�S�{a��9y��d�l�\j�Ϸ蠆(/�{�-��ذ.�I)ہD�B�G��P\ɥD�ʹ���Y��m�.��N��T�����_�ト�_���W�V0�O?Z��v!?��{R|v�!	ΰ��Y�p�0�k ϼu��c�Y\�HI�����	�/⽒��m�E��4�ў�v@d~m�C/uvd��}2��$�ox� su4�"*5���~D[fRe�Q���n`��!k��Ҝ�0վiBȆ'����Z|ŔM&]�I��BJ(��4���]}�s��YA+����� W�Ԟ�ġ���Hr"|�9 �s!M�gD�BE|BO�]�(@�Ԑ��g��Lm^y��4�2�i`[�Dh�g����Tɞj�2�VVN�3Np����]	��$��I/ ���)z�l/���v���K~)�A��/�JkάB��E��n��1�sHb�uZ�&��\h�vנdC�0����ГRA����vk�djZx��,~�2���5p1�Cyc��Lo6*����O�V9A`�QQ�������I�ϥVɦ�n�Mu�ͺHni톧���B2��#���A�5� _�5��]U`�^���2�(�o{=+��3�2狗rPү]+D�0������_v��RQ�Q����-��`�b0����G'��l��(�
��w[EU�Q~�FUvk���ܖ)h���i@7+�ь��	X����J�S�处XGCI���=)�2<�����R|������Q]w��Z�=fZu����4�:ߺ���J��:� ���yd{�r9�v��kc5wz��?�s�%x��;jW����\vJ=�LZ��i�b���'�s���LnzOs�?W�mQ1������>B�`~ԌRKg�L�y�ָ6�7<Wi
�����7(��DAK���%�"���}�7�c�\Ƥ��� �<A�<�c���A�������^��h��ŷG��!s���F�7Et�0���m���W���n6��s����'e�OĽϬ2ڵ�$h�Jg�`�;�%=w�W���MuD������}ef#�=O�o���"����:?�����+,�����)&#?�`5��
?�m��&��d��������c���j�zbHv3C�޻��7n�����u^e��I�罔J�L[�:O�ڴW�,��b�Bɝ����{Fd߹x��6L�g��,�'����^�1�9u3Q�^ܮ�&��x�MU��A	����a�\u G�"&���z���A�l�"¸w6�h���y��_����,PJCM3����k��%������Ļ���L�����|"P]��f2��P���Y�t�6Cz&l$�?�ԤV��]4����K��O=*�'�L+��A�2�rr@�-�_�-c�l�e8I�k��%h70㲳�7��DBМڤ�ew�m�1J˻��oV��f�H��ߴ�}���M"��|.��ڦ�߽�����ο��v�>������@�����Gm�WbM�������^��щ��إ�o�c��'<aX����F!�P�L�-WG���O�M��&�{�G��电����·�Jv�z��T9+�^�acN��ʿ�W|o�.�qv6:�|廄��B��,֍&��R�M�N��%P¯�����m�lW�i���f���ΛOM Ox�M@�)#��ye����Z����`v.��*=r�'L��$y�N�9��_��˃�u��"%c,�s������H��>�c���1��`@D1�J�,\Ϊ��5��+��Cb�? у���õ����I����Z��F���M���n3*�z�����eZ�&Z-8N�x�hj�-��~�R����aA���l,�8���۴P��?%��k�PJ,�'|�U ��$'MT�7�-�La:�f=��HQQCʺ��ɂA�B��FI�����Mb*h������A��c�<�JX6�����o��'��+z5����Y洐.�+���!��-L�D�(�D���.�����i����3���8�)�8;CNB9$�ޅk�K@��yϤH�i��Y���`���d�(�fƖ�3ǚ9��My!���(u*Wy�ŠBQ5Ks�/����R%+�!��{s�i9�)�"�,{.�Z3��@m��
����,�����n�J�`�1kPE�Dg㆒6�@�@WKExm���P�[X��^4�_�=��
R��R�?֋B/����`�e䰤�b3��(�c��nJN�����nQ�Wp>�����!��t�}D��eҤ�q�<�^��T&B&.F��N�\1�g�U��;���$N|��0f���bѩ&V��ǵ�2ѻ
ʼM�]���0	*W�\w��϶����)��M��3�X���{�Z�Z�]SW+�b6���34��QEX�_����Q?ZWWcז:c`�~�i�[����T���Ԅ��2�R� ݉� *^����O}JrE�SC��N�Y6����t��2�\����׺�4ߤ�����Y��X�"���^O�
|5�zv�:�4��Q>�-�9(GA��k>�H
K_g����>2otS��<��<��;��]���ɢm\�F��6��ʨּS��e�M��%7���٦T	�y���*�3�䁀?Y	p�`����ڵ��IIk٘ӝ���4��ې��F7m�pH�+�g��j�W�c)������R�P`9�J<	�.���&�k�~�@����j��4L���W�	F���3�����%�6�|��z?��_.m����zYJ���9���=���(14A�^�w��\�u�ܙǯMs^�#ƙ��}Wq�m/�������^���N/��o'eS�,#s��>sТ����y�Sz�9'~-w#"����o�aY��Q�s�R�:��,=�B�e�x��ʞ<Հ~���Q��ۂ!AC����w6�G�nG����`��Vm��|$cR�<�蛵��`5�.~�ď���uCq�w���{�Դ�5J��߸-���ݬ+ޟ9��|��?�tO�;��ǻä4���`{Y��"8f�)!ٕ����(�,������?r�+�Hh%����(N�_^,SXZ7r����o�l\ƔԌt�p�2��3��o��6����R�u��n'@lǇ�Ɇ<�g�~h�r��߁2���U++Iz���װ|�:����r����|IS��<��?n�c��ʟ��H�t�����{�z��(>�Q��+-�5�/ߐ����*L?��s��faƁ�Po�l,�X|B��ξ>�H͟KWw%��Bg��#o�P�����y�:�jb�fY�-�b����M�>g�viN�9��$t̳�<xˢ�/�e�� �\�'c[��Bm�\+~3z���G���ɣ6��Sj@܅�x�o G�=&2��Tѝ͊^2��x�p溡z����lGhR��{��b)���z�����]�X��k�ZG'$d�Lm@���ٶ�t��A6��/���g-qm�g�8{k�t�#�h#����5�&1���^�~��� ��b�+��� DyJbFQa�,{�`��9��TF��F�����C����=a,��̘�.iަ�/ua����W
�2덕�J����d8�L��S�G-r~����[��DW �	R�:��l}AtȲ���~uUl\�7�pD���� �w�l�8�8ę�x]�М^��7u5��ṰX��{�į��ʣ5#�p� �tRM�|bK�'�IH�o�՝aη�=q��'�9[���1ޑ�茣xy���wb��04�W>��g��TN/���Ql�|�C٠�7B��?V4آ��?TߎԆDSX�PT�fcǀ�/�N���y�ts���G��:�Se*�%��.o4�~?���Ch���8b�;���mɞH�����=��?�u��^~�H�SY �+��Ֆ �<h�>8^���?��n7V>�eg̟�I�~��Lʒh.&e�_ �����?/M�~�X����"�s.Vǉ�@�mZH� �*�p�X��@�U_�O�7�hYW���#6��K�S]�>�l��h| ^a�?8��3�%]L��}�f���]ⴗj��H=g�{�U�I@��m��zW��ka+���@$ ��I�'�K�=�-��22T�� ������	����hwE��{� `�g���̠S�{�*��R���r�ˆ
3߬]�gK���9��\(׬�Ч}�!wY�_��'j�#�u@���i�Y��
�@�N �$����\F9�{[ɤ���i�#�f�bF	Z/mOP O���r�drѯ)���+K��� ��I��L1u.�?V���;�ȿ�Z���P:쫄���FO�o%G� ��j-�ʶ��JݑA��:�Ba���!u�ʍ_�\�Q�˪KP�3?hzM�7e�&Y~�Yۍ��hc�o|�7���E��oN%Էk�9jH����X�	'3j-���b�d�`a��ӮW[}������	I��S�"�+�3%�x �M��3�,�#�Bbr_��D��Q�l6�5���e�X:W�/alU5���soQ�׽�eޙ�����ݤK���\��#���J���%��z�Y�M����Z�ū�0�
3-	�
=���z�<�ȸ`��gPZ�0��;)�%�6��7�ώv�
��q��D8vM%�c3���~��KW;jl���3�v����|ӳ�
IDv�}���TDE���;���
0`���t;JrE�ϔ��HT3�Am��B��{�R���thm���Z��1	�eo����)/��5���?��ϕ��O_Aol� ��<T�#Ԇ�����{_(pH���i�4�ޱS�N���+4N�]IJ�I>>�7O���͂d8X�S��B�a��a����7XK�ц��!kB�U��@�V�N��h��j�y���C�u�ՠ:A�5�ʄ8	�YMW�� o"^�<���t_	��8���2�L���0�
���6?�:Q��~i
-�d'��f�a���	�)"NɥTA��OԘӔ�j|o����ޣ.���e�CN�����܉O���%3kt��!����0�o��e�%o=�W�
A�f��~G�|��]�X�@��4����P�͈(_q���һܖ���w������y�km3c�C���_�H�t�W=����}@��Y�goC�v׼�i��G�_+���\O��([]�T�5,���r�mI�J+����\D���qͲ9�1�����
���!���L�j�r�S6P�ѡ��p^���k�J��7��R?ľ�p�����0"1�7
��>q>�&�͆�i�h�B���?`��K{Jƅ�5��;����Ph&B���L��/���;�~|��-���ǜíV<���O�Ap�W�'�:ڹ���۳z�pxҋ�ƃ��	)�W�e�5�u�u(�p�Zx�������l
�_
gϫ��1�^�űѳ���BF⿒�̻3��A�|}��jCl��䨏�(|$���UY���ӽ��r�s��?�ohe�yp�Hq-���_:�nz0% >��� fk�7�x�������4���r��'b�����ɾk�t�r�6y���W���&�1)�P�:���� �/3��_ˈ��³�T�q}1��g�I0��-oL_��z��-�rJ�|�����<�3uD��h��_Ҽ��/R#8C��C������3{l��R�lK~�_J
\�&�A������~����n곚���������b���v,#׏-)�x�X���~:����a@,jF/\ l��V���3��cſ"oȎ$��M�z�N��yI^fmX_�}u�h�II8�Нa��a�O~��t1��ؙ��$�j�&�J�����죡�pUbC칧�-,�VntMKL�#;��]5>s����<��x�ZG��Aֿ��mBch��s�%�����2��������j�!�����<�4S[X�6]�F���ߛL��?�F�W���(Y["�(�
����$��V�w�zl]y�3���Ng;@c��N������9��3n��sW�/İ�.���'P��|dt�͸8�+n������u_o�g!�K6��6a��7X�oMl�;p���7��e�a���]
#3ͼ�.�Qb�|��^���R?0?�G�ҳ�S#w���I��5�H��)��o~׾/:�g�\�a_�RW��&U�����7繒p�p�
�Z�͂r��pxZ�%i�Os��3wv%A+%K1	_G�"��\���Ǝ�.�=z������ �g�8B�Q^�`��/�r0l�@h��w�POm�GڗRa�J�pY�`T��m������>6�[�G����^p�MDB½V��U��hY�k����`]�w4*���K��eC�Q�8)�W������v7��He�I�ԅs!!^�΀�?�_&�>&XU�+; �h=r�F2����#+��dU ]5Y_u枩��JD颏������Ӣ%���������wا;�j��
 �|���{���B�̮:����k%�����1L,��4F	�呬�	4������c�1Z��
c0s����v�Ē߫h�a��*�#ʮ.g׿�������ȥP��[[��IНŊ;p_W���r/ї�k�L��)�˨<A�����9\b��=�[�Xe�b����>�]�F�J�$��9�=Ԙ���:B��q"�ը�'>�)d����u3튴� �i�]Y���g�A=z�OuB�7���-j���Bd��ĨQ���21�⿞>ieڞ]O� ����қ�䘽��g>W�|�db#
yM@�|0F�nE�"�O�-�)֮7��X�{�5V�Y�j 	�$���Q��.k
� ��K�r՜ �@+���6`�Dg�8㞷�\&�Zi�Q����,����!_6�=�i�פ�p0����e�P��w�'B:n@n���m�������i� ��uqoǵxM|=�:
���0�����llR��+SG�;^Ɖ��7���*ΰ�%�$�/m��F�2�`If37 �"��fI�q(��8Z�:ЉRml7�S���
i��ô�
���6Ck5?�����jmI�	�6����YwP{����W��ǟ3�q�k
��r���7�Q�S��c�1_�Mk�)Hy2���߉�`���ⳋ�I��=��ڗ��e�@��NCܿ�������>7:�i�ey��D:+���˖&c%fX�o�Ԩr!0�v,����J����g�=����"8�ʅ�(��Ϸ�K���V�\-�rP�^5R4�Ԧ/녟����\�6��O�p�!��č!:�:�|V4qx�Y*�uQ���7�W��H��8�Bu?��e`k��(f���/2x)�5
��ɯS��-�_�jm��i��Z��`8-+"��9�|*�^�o;�uY�RnH���KN��� "0f�w��Bs�oA@��ḷ��Zc�k�L �n� E��N���2�:�ru�B��jE����� ;���=Zp��M����QF2X�9]��Ӣ�Cp�\F��/�v�v��=���<F���>'��Q����S,n�<f�C�1\P`}MU�Ͻ�`�r١+�*5�ktw� �,��,�X���ykp��F�韒#F�c����4���A
�5jW��<rIb�W��ꅱW�[R	NZΘ���}�"�]�\�g:ۍ��~�{�HoQ��Tk�V�珀n�1��=]?O<�\0NÑ��7�u��xT��I��Z�t��֚�d �~S�>�uH��+����b�$ױ{�#�J�63�o�D�A���_��zʀW]���p�ԝ�
%��������e��h�S l~�IN�e�!��kqD�DG"3	[ ���y�Ƭ��2'i�� x^'�`��9�oi;��+��Ee>��M�䝑~�:��c���Lm����X�d˒�E��T ���8��b��C�q�hC������%�N-���ƾ���d�{#���K=c�y�����T�d͍H��6 #�zis��m�G���NA�^6��oأq~wؾ�Ys�U�ze�?��3@IJ��l�m���Qm��֎JZ9pX}�.��ť�e*��&��|�����P���:�fGn��I��'�R�rV��~Nz����<{6FB��U��4N;�s�~%�t�p��\ˤ$�X(�}��|g��~�a㚇��E��M���	��wkZ���bF�+��y77,]�XV����O*�l�zQN�zb���{��.�nS^&:A�G+�i�����y��MΞ\�F�2���'�F�n0�@:�1��Z����J�S�.��/�Q!E�I .�g�ƫ!��rz\��U�a�,"�+Q�i$h>�Sӏ��7�o[�D���[м�W^�[.�������r���!�����Js��t?��Hr-2���#��f�AHl�0�Pw��l�d��V\�um�;���߱�zY�s��5���}y���6�=	�B�$�-!���ٿ�������7t��+uĔ�$i�o�61K�k��$d������`�I�����E�ƪ�[���р/��֏H(Y���J1\���g^오6�b�+R�.���A�ۢ%�����oJ��F	С�j��Q��q�$w����=��H�9=�Z��P<��h	��CH|y�"���x�4�YxQ�u��]hn�|m'	�y�� '��	xԵ�E���桨�,$�aS�S�\t�$��%�iӵ��m,Q`��Ͼ��iODܿ���Z��<(dШԂ���j,�R@9��3L���\Xh@���)��&�Z)�g��-��qp-�����j�AY΋�;ѡ�`������@ae ��!O3�ۦcT��^��O�w�(�^� 5�_����dQG�u�"jW%�H�	��a8)����k�i׻J\�>$�Q����|��&f����P��v8�|N4�$8���~���M�[��g�$�Q Wk��*�UA=z=w���"iE!��YZR ���{*���ŧi9��V�z{g�f�A�C&e���}�B�������>��U/���s��#�����
�A
ԑ��'�1�LG��S��CP��od-�5!���,���� ��z�����b�e���l�\�[S�Z��=�e�it�a#����1�cĨc����v�y��J�"^d��~��4q����̂�!����&0�{���"���G���*h�H���?��˺� �I�ۢ��&�]���s��Fx��m�u���Tv���oV��Zmې㤘�cxw��.abJ��dd�#9:0��2)������Z�	��,�PSᛇq���/��p��3�:�y� Wf���(���ٚ(�K�ZM���sK�L�eFĿ�N
�}%�Q^r�̅�:����vg�I�R���"S���f�^	[?�_26LR�|w�[~�ak�.����,�޵G�QQy�3b�'�Iע�� s:�Mɣ���$#��JEm�=`���v��tw��3��t�&��g��đ�R�yj�ڛCK��ۏU� ��n3X��>���ļ�R�๵���g���k?�y+���s�Ǉ p��T�n�pY�{�=<1%��E����T�WX���>+�"�D��#�B9�oL�_�� v��7S�I7�9O1���0o�~e�h�8�m�n��. ����<-��'�������u'�8�J�AN�+�:�Y��,������ w�؃�.y�H�a-p/^��L|/ ���Rʡ˞ :i�S����(���"kX�����@f�����t���J�nb����U/���MsdF�x`��՘,�!
��4��1�g���L�e�j`���s׽��ĵ(��;�@C�K�P/�>����j�AK�e�����Ҧ�K�Ko�U*/�P���
��B��%H@�jj2�M=j��Am3!�A\o�]�*��������h���l��� �؟T��� ����Y��o�+��I@t��68�RD�P���
Z�=G��6��=�y3���H�*��T���xH������6���Bᓋ̕(�ۅK$L6��툈4����c�BbcN����[|	F��1ڌް�	d�g0�]Yx��yNC�s�n�H����]�uZ�����Z�#���L�{rq<qO��6�`��wa�`�c�v�G!�R�,/|T`D��S)�T{�M�^���{�ʘ>�n��Q�-_��2�81���<�l�~0�I?y��px6-tb�y>5V"�ٹ�� ��8$`����"GT�B>�}(��o�W�I.��f�y��a
ҢgV�p�W����+6�އ~$Wk�YƱ2�K$�N�5���'�z�2���c�k��,��&�v��(E��[+�'�on'm`G��p�"Fj�!B��3���Fln~�&�Wȝ���@��>F��ֈ���Ƹ�{G?iҒ�/+9���>܌e�w���w�7���uc>���@\[e�z��/���Έ�O�5�	!U@h�(��a��PQ��J���A	�G��i�.����XF6���#�厱����]���V������~ق�;��
� ģ_O~���T�L��x��6KU�E2xY��)E�LU��r�^��3��3��D�0�`��M��	m�jh�-s.�w����+�`�[����&D���xH,�,K�6�M>���\�'O�����{`���	͕
V}9'J<ᄺ����
��z@�g4@�p(Tg��R)�Q���ǿr�a�ו-����p>��XA3y��=Ҹ�gl��t! ��p��$ Y���lM3D�r�_
�7���̽��/nXKh�y�͸�4E��A�c/o!�Pl�ͫ����li/��`}2��'i�܎y?7)*����'�"�B��Sf��o��1O��~63��3��)Q P-C�q���OR)`�IAǌ�gM�a��@<�[Qn�(D�o��Dݾ(��f
�*v�ܯ�JTx׽U�0B����瑹)�T�x��{��
�Hcf��Yx�N��T�R�S�r& wn�K;��Vx��q7���G�ux5��}8���E�G` Be���G�wZM�#����;��\�و,����8���j*aB�\�/�9�QLk�����31�_�\�crJ�1�����;����=ʊ58�����[O����K/ӟ�����Q���I,cb��A@���?{b|��/m(>�� �]���G4\:�F����R�t%r�,]r�R=�|Ffñ�H��p��$m6�8R�����"�i�V�W��fI��pJ;78�3V�t �v�I��6N���*.�=x���Y-F�:��S���i��ŕ��*|�w��Zgj棌��I�m�U��m������a:jɒ�:N��so�&��`��t��Kv��d$����.����)�аc�U�F(�+qԋ�I�#�YOg�����^�,�$);���E���nDiU�u>R>ź
7�0W"�Q��b��A�Y�{[��y�zFy��e��t  �90�v���%
2�	���=�/xl��#:���u�*���P2f��YBa_�cAB�d�Q� f�w,��=k}����Bڜ6=4��d�w���v.���&(���^��������sy���ѓC���:^#v�;���ɧ@�M})��;c�dR^����!�@ۊT�9��8��3�b��o(�%�K�G����)cW�
K3����4����[ֻ�O��^��B��r97�#�	z�`!�]Zgƍ�?P�B��:�.���.9v���c=�M[;�ɣp��gCr��}���L*?km��� �,
ioK���H�����p����&�.�M=ό��١��ymL��RDn���K�e�  ��dk�K�ʚ1�_q*ңn�r�]��A>��_[� ��9���h��+F;���xlkgY�h���Z�]%V�+?$�"iӭ�U�U~&|5Hj�py��X5�|�P��m穈�����
Y�0p�=ʠf����[=���@�Ǵ�SQ>�@w����P=�"{��
i�u�*�y�/N��� �k6����bs�ׁK�]?e�XY�呑+�z��-Y��["���m��ńN�l���r�JЊI���ѱN�*{r���&=x=|��QMP.��y�[3:;�ÿ���g+��1�UF�1M�z��{s�$�;�g�Uq���K� �͖�s���͊9+����sYmD��ٷ+b�D��D5��s�%��l��e��q�����	������CbM���W6y�^�^�A/��{({�[u3�}��/')���2��j�feB��h��]���C��`aI��T����n�MNަ�.��q��΁/�&u���jG���,'t���O�>M,㍗;cU�j	�σ䛏 ���j|���Ķ����U���K��}��� ��ٗ� nx�7��ˎV�=H�ͩZ�	ym=+pK������r���Ӳ��<����$��T�	0�S&�o�{,�~/�h�oo\ ��*Ta�n��¡=�H���T>8Ӳ��)�L���T�i9x[L��?वy�eJ����⤦@9x�ߎ�ckj�H�ZmG/�|�FOo�#|W�\�N� Y���Z(�x��V�Y����a
���!��̱�5��EL��<
B���B�X�|{O�+-�^=B�f��g`�tH!D�o���Ӓa��e�����b�"�]��h8��Be��V�Jh�i�Z�� =Ӕ�Gk�h�E�0ȡ#�Tv�d�E�u�"ԭT$,�yA��#��er�2=�Is X��Ҕ�(�KA�_�%]��]7�{�}����6� �J����Cr|�T	5��_ђJ
7�|�֗��rǆ�7��dfcc��OtV C'Ye�}�h�T^3�9j�e�5L�R&�M)Y��5O"X��m�)��B�0��O�U�>龓_����F���GN0�>!-��¥�d���Xp�KI�!uW.���9��!�]O�����^u>чt��2L/܅����t�����z2�c
w�.^�fC�Ux똴��(ɰ��>�D4L�������1䛘�b����e8bI��z�*��.Z�Ft����g@V��9�Lv99��qc^�n���@(��A�(�%�l5Mk-۱�-��1 ���F��ܢ ��%+�Z,��hzQX�0'݉�<�Z�$�:;��@����kc��>��҂�q��rᄩ౯��vjn|]**���.�(]�Kd�m+��+}�k�K���n�Y�׉�[]M�J@��<��^q���c���a��#z�x��~���g!�v�5q���ʝG3�kX���PIAћZ��R�-�GSU?�9,���'�����vV���?s)�>�Z��?�������ۋz	����TQ��}p����wQ1U)c��QB��-l�8$U�3�1�M�
��xt�c��YK��<��<�1�A&�3'3LM��W=��N�v͞���E�]�F̀:\�VU�w$)�>Z��R��<=�,ݟ>r��I��sm��L��r:�lwۦ?�r����C��14��H%�(���lz��t{4*8wU��./N��Ϋ"G��>D�d�^�����`�18��1�x&�E�������ͷ�`��f���$Z}/8��N��fcP�/���R��c��� Q:Xp����~V��Mgj�}� ȳzSן�&N#>,?���#�%H�֌y0�W�ɾ#L�iM|N\*W�3�~Q�7�����#l��TM�@���w�GF]�u�XWs���7�Kώd����h���N2j��B�p��dm@�G^��UE�^R�>�,jU�����3�����Ԧ�O�M;�4@��vؒ��i,��7�%o�D�@:*˳KQ�Lw�=���� ь�z���	iד0n�{$�����?tg��ڦ����cBAKa��X8kW<h��"�uS ��cȏ��;[p*h�ᷤ~��|}�-%�L�]Ĕ�ꃻ4��{����.�#8���k��-�BZ��CĎ�6�pm��-E�R�g��!kTЈ��Ȅ΅�a�A�A�����j22��oxP��e�v)O��/��y���'m렞Q|��
���+B��)\�*H>ퟣh�?t3��lx;�b�nUOr���Ԭ����_i����B-@8Qʹ.��{���*t$�νW��n$n��zq��:�t/|�,��2�R�=��E�;�����01	����t��f�ER�}	�<�tPT%z���h�q#��"�ӿ=�@_ ��qZ99�N���T�4�(���rށ���G-�Z��<�]�A�=�� ǳ(��ܥ��yPWk�8]=���@�9����>�#��0볞��>E@?~�(�ߟa��_�?`&1�!D�4��<�D�|p���9���)�"�C�Pc�4/e��G�=�z�e���-Q�k2q9�?\l�����˞h<�;���c%]�ۓ`b������.11�]��KQ�g�]�a�q\n=��h��º�~;fW;:�tYpg�v7(\�VȲ߿j!)*TM���Z��@a�QO38q�4rGQ1�� ���R�'8���.�ڒнW��2C�2j>����2�U>�W��y$��Π>'����<���v ��aG��c���lߔ�8���X�׎�Ͱ���n� ���8#��/�>��,���u��{W�t�C�;�5� �Ԓq=�Og�):�o�,�UX-Q��
訶 ��&C9)�3j��HU�Cn	�؁>԰��!������rΔ�l�ì^\1 G�tk��v��( �<f�w��kƶ��������ُ�����\f5����鷕���g�7}x���0�5b4�4ꩅp��iV����/B?�%��"ף�>(-� ��
���l���k4���u���μ:eC���������W%���r���"������F��+��®�/�������=��n��|}���6�05H�*#9�<� �N]��	�kB\LS4UZTK��{��Jo����kn����U�<PP5M�}��8t���~��$AO*Y�k�TL3uG]�]�}#r1.�4��;����
�;�H-fɀ��P���~ׁ��,ś�P�!*��t�t	��h\�Z����A҇� �C$8�J3�]�zfX��F������KBl�!�������1Ո���ZK0�Q�ʨPq�nFn#���;e9�Du�蘪��������K������ñu	���%e"��.a�G���Ca:N�	�L>ݒ��s�����yt�ĲP%o����Q�>�a��_ǒ�4�L��ڍV�D�so;(Ŷ$�b���k�c5O�����Шa��?Q�����n��F���0����5�I�����-Gr
����u��R�b��<�#�@�����3@&I�d���U�����9���w�&�/t�EA6�T3L�Þ�0��@��<~*�k�ɳ/�{p6GrI\�Ía!Y�`����=[��ȑ����@���/u�[�ھk	*I:�Ii~ H����T���IBQ�Y�Z���32�v�a���̳"p����8���melVօ;ҋȪ1ʴ�\p���r_]���J��"�Y9�\N��~��\�0a;Ӥ_�q��R.+W�1O��Z��x�g�1��Y�9����&��x�hg�g����a2�#�n�̿��j��Z+_����m�\Y�.}�9j���퇐�uL�����F�/!�\�,��!d��t��|"�ö����ye�>�Uլt��xt��L'�=����� W\�����'okn*)��J.���1�8�G�����K�t@-7�f�s ����:���
I
�I#���U��
}&�Z�#
<�D�G�����kJ�Rڭ��|�D��<��K����-��OW*�,�șa�G��R�h��oܿ' ��rhb�%P�˚�=�Z�Q���F�	(&��cJ<�d�M���,�n�=�B�{�:9�WEє�44F��k�'�I� =�0���bq0�"鬫K�e���bm:=O�YigT6z[�Y���G��\�n�fr�,�$����a�Yz�IE���x<��}��⿼m'�^4�qEn�ZB_xY��.� 7&� S�K^�<��d�{4�ԧ��ޠ�?k�F �I�#�בӉg��.��'z%uX={�G�H��dD��U;G8J��M��҉gf���|���;�)Tq��>ـ�$b�Ӈ}���0i��z_N�ͷ=�����d�v�I����W��"�|x���=�@j��ArGaܗT�L�Kq+��ے���k��e����h=P7"K)s����_'���'�H��C�Br ;bZ����P�+�b���Y��KBLs���liw�B�����y�B���m~a��=:"dl���&HV�]~R�.���W˧�U5�����&�\<��E�����2�"}��jΊ�R޶v�~�H(G����h��L�v>�/�U�� 1�f��Ӌ)��l(vGl���>����.O5��]��j�1tyPd���>�Ft��nEW/��J����L������U���~v��:8��@J�U<l��[ڀ��2�Ǧ����f���݌���1-5)$�����)J\J,�B>���م��>�Չzu��XLr�<T����(�`�:zrk��#N�,��H�dAG��2\����`�������!�H��,��hK��}OU$L�Z�?�����|F
>�d���ް�Lמ^|2�4v�������k����g2��n~W���L8t&�?���j��@���-��
�n8���p�2,@�F$D�Gj
�,�H%jz�~RkH\� �6gsQB#�����ud��̦9{�D �;� �ª%��,�O�ZW�i�	S� �+�N��T05�yۗ�*���R��V<(:�a�=#�l�z�P���u��"�g_�� %��"pX���k����,6�4�^��9q.jY���8F����"0+<�Q�^	-�
$2	����������瀣�`%x�!~���m@x�r �������A%�hC�x��n	�^�'���pX��A����AtV�ӗ��A��Uw��@�@��8���SS���#�]!N�9h�o ��6���F�K$<,l�E$R/j�K~���?�/��-Ā���"gؿ��Wd=�V���d>l�I�)��G�X�ﰱơ����wF��&�u&Z��!E��� :�B�.��#	�����ሄ���'@�(|kF6�;Y��1�3C��J)�~�n�T���^h���ҵ�Xw�����!cF;e��
��"���j�/m��r��aQ+!�<n|�}�����Y*Z����3s�����֘�Z�����~.��k��8$�ޔj�/2�Ӽ�*'݅�[�#��߷�,j�݄�Ф����ks��P�����נK�h_� �}�*�+��e���V����a"�4�6*�2S�>����_\�����a����.:�y���vI����Eo:l����X
s��
�+#���I�h�)s�[3sI�YS>k���^�8�,>l��=�aL[�� 2
5�?��'	%��b��L������+�79-������g����ְ7n��]S�u9ky�i^,h����Ŵ���{��� ̅�0a*yS������cH�ā$w��NK����ʐP�٩�|��y�Dux���S'S��d�v�G�.F�&��Lˇ�ܩ�ַ�2U_�2L��,��L�����zz���S��P���A/�-���PqG��LI�<�Z��==`�
�C�%g��4)RJE��sU��C$�k��W�%[�7�(:щQ��h��^pÔD�g|�]�p�Q��j����}�:��C�e�,����	w��Q�JVooN\yϓ��X#N᠞�',ؖO������+��;*a����?����	�R���N&� <AEK�)�X�	F���Z�k�Fj)��w��a��i���P,���=���fL��WÒ+��C^d]i��ڔ۳C�)$b��Dfv1�|$S]&�u{��y�N�3�E.j��֓I�F+�xK��V�r�cC V�O�E����C����R� e��!�,���C�s���a�׾����Aj�V�l7�Y�W��e��N0�-�,��9�E��B�W]lWI�`�j��ѠN���#]Dr���5�0!�	r���8,:��(ئ� 
s':x�R�?�I����F-��
 �A.��y�%v�d�e���y��$k	����1ݰm�P0���[|�ǹ�@�!T���J�7�����ȷ�j���C+bw#:P����MM�C��U�m�*�YI£�����L��Mj��P,�_���Ն4�Fw���Ҕ�:b ��&@հ�R���k4�v�͖zGկ?n!ܢ�"�4�w��f�#��[�t,[�k�}�{ֵ1yIu?g���E����P�(�S"|�_zq�8R�K}�I���.�X��n�Va�HoY��ώ]u��u�,E!\�n�ё��Nd���D���b.0Q��L�~pR�=�^�9��݅�	�(���<�]��BA�����%���<,����v� ��Z����=�~ e@���'��Tg�N$7(?ȿ��aZ}`��庚~&�)w�+��)e�#J�����h�-n�r��v�
iC�X��o�!��=:�7��V�M�0���*~i�j����B�b�Ͷč�EF���oB'�+�[:�^!���$mF��WwÑDl�4�I��?�>h��y��(Sm��a<	1������Co-i��<��{s}٪��夸<�\a�2�K�W+D���!l�t��`׿��w��r���W�����+�~�F{5u��#�o�gQ򱼉w�-)d�m#��y6��{�P���&��7K���z�M�����V1�WRѧ��Ｖ'��4����J"6*dA�4���3ס%J������~�2\��e��OK鼠]�@���J/N�
t$�}�5�H�>�2��= ��m=|��M�y�_3&�:E�����i��a�ƣ�?~C��,�?�	�P�	7*��YW�㥅$>Χ�:m�j�5���a�@���a�jY��E��uJ��?�ɋ�{ى�U�U�3mEo˒�l�8�AM���:�"�6���%%[en�����$+V����7>�k���X��p �-�a�q�;ph��k�1��[�{P�J$r��P���?YbJ��?)�̽ ��@����uX7&8ׂ;Cs�X��tS4iO�л�C>��2�G6�:���gyp$��>f��*)��p�e�ﺅV�vV�S*���� ��=_�E��$��C�مL+�W�w��J+��W@,A[�D���3	��7����{Kbu����%M��=�q����.ؓ���}������m�Q/���Z:����o2i��}ZF�<g�묠��o�C����rz�ď1Lޠ���6S5 @�n�N���<��r��Cu>�.�c�U��VZC:�j�Y��+��զ����#K�-Q�Gҧg� ��Ǌ�;̚�9ǛfB�j��dCXVD43ϒ��~(��N�i�lM��ʪP�;�M5�6v[�y=b>���_�b2�+�y�vr���,���d�ٽ�����:#/�q]6,0���+�k'>J�.�ęn�o��Ϫ�H<B�"Z>waO����]�cp@����V#Z�U{K3��L}��U�7=>-5m���ƣ��P7��� �����l�N[�ۜ�O��b��A=�����ud2�N�����qFp�EF�K�v��A���Q*qe�ҭ�d���&���OFMFJ�#X�66)�����ҤҸ=TM�e���)��>��,W�����F���ð��:���Ľ��)�עayQb���?q��)���H�2]k�4�E�)Wx�R�[�*I�n�\T2 ��.B���KQ�4�ڀ������׭چMF��``����E�p�ҪƳ�?M��)n��|_�16ޭc�|�:��*4����n-��Һȭ���v�_��[
�g���3-u����K����������xl��/�}i ��ޚ��J�b-y�1(�#��<KD�J�����V���`���~E*��n�4�]�e���2$������(��K�ԡE�b+�bpAa��D~9々����}Q�`A�1fO�jz�6�l�'S	EX�a{&6����u3Zn^�R��c}��bGޠ*��Ż��i0Š��~��7Bϲ�?9Ӈ��$wvs���f5�b�i#��
�d�2w�c�fJ1uG���]��"�]3���L�/ѽ��)��++K�.�ud	Td��&�6��t4�=ފJ��*�!ޑs%�<JVb�����4!�����-QRK����Vn��M�g�)��1�0�e��
Ab%���CD^��4#8�Ld��� #�ɟh����	�kr�����٦+�����@9d8Ip�0����4π���K���	�[<�O�%���S5R�W��8�*C�|M��w떮lI4����z=C���	]}jP�P1��۹A����� �[޷OO����`G/��큢x�s����`O܂�(>�$��+�x�l�YӨ~�L(�ʄ�%�"���P�#J|�6�o�?z������%4e��FR��a���LQD�0M�.l� $���6�r�E=�u ߪ�k��{<>7L��Ě�)H_f,ˀ�4����=��۫GYDA��\��,e�I��]
��Q��T�-{�M����e�� �gz[�.�S�C�Q��k�7���WY�2E�l��7W.`�Y��c^�]��w�e*v��<�#��@��E���Uz�A�gֹ��,�Čũ�'$�b�����_A���đ*�q��=&�e�����f��Կ�E����p�	��d2�)�<ARR1���Z�6b=ܠ���k��� 䅕�ϻi�Y.��q�Z��"�\1iF�˹G�mW�X��`L�:O�GÓC�J�=�r�J"���|�k���w�dwl�\S��-����}`�6��M�Kƨ��*�Ky �����kQ	`[���z��g2�åbkƸbk)^�X�_�7�Nyo���Ϣ/�)��H-F��U�3�Gb�(
䕵\�@z�z�,��݀���
1x���-j l������`�3���n�4
H�8�M�]nT��Bf:��TL�nL/݋Rv�W#�8�vfb����?�W8+����:|N:Zz�1���I�����Q���].�����8;�F��T��tc��xSflXk��]���ʗ�䈊��O�%����J:Rfp- ���K�"3��Ց�{Jn:��4���N�(��zD��U�v��q@��4��<�,`v����Eq�r��e�E(&�qZ�]��?�Ng~�;��=`<
�n�܇qhZ���������f�5A���b:��L}��8�Q��]��[�&x�ꊡa�xzfe��w�����F�����-1�k^\>T�8� R��o��>�O0���J�?��1c��]*c��a1΢��;��7c��2v|
[[$A_����������d���kԃI5���,󉠅}�S"L9�,�w�궥r�`5��E�wYC�J
�bD�	}���aZy��ΐ��ͥ��M���cXm�'��ܘ��5c�v~���/�h> �i�6/�x�o**�j5��د)ِV��MI��05������ԯLl��dR��2�eTe<�(��z���{k�� ���P�r0�4Ӌ�bLqDa��G��K���ޱq�0�x�9V��'���u�F���yϣA$���K�QH�)۸��`���ZX/e��׋��j�\v�-��s�݇��:��]e���vh���G�T���P. z�&YN�����bf�''�澇4�\�޵1j[y�0+k�o��N���sI�垐���=l�9�	Ck�FZѧ�5�.�I��O»��û�%���%;���*�����i�񞙖g?5W	jE#�!ő֧����c����wķ���N�rv������"H7�tB	P��4Ty
?��q�6a�A��Qѿ��9)���B���~�6����{����.Z��n�7��C���F����=�n�ʨ��2U_o��y���j�7�Ԇh��xLT����09$^~��(7�|��t֦ໟ��_��M���&�F�T��Ҩ����X18����BtFP�s��`^3I�ƄO�iC���������^������oz����n���j�NEj�̒����Z���X��M�F%Ez�}k?ز��j�����):o�&"g�h��TF���ԣ�b�:C���:5�bK#���@	-����|>:*�%�c�HY������OH��y	���pL]��{��"�A�3O/�q��p^a�DH�h�}�����(݁R]�>9�F�r�j}.*hrv`QN�E}sKH��E��ҙj��ѲB���bHj���$@��qFt8R$y���!�&ؖfJa��{~�
�i9���[��}g���6�c�6N�^녣
P��xɕ��6�г&N�ӣ��waAQ�s�tw�OL�q[x7R��8�w�@���8������V�����r�.�}��ҋ�2��]��_&� Wn�C[�	�'mƀ����V}?�%�!fY���n�(��+�S��v�n>p�/�"�^RPP�D,v��at���`���]�^/q6bR��ɨ�%��;�$P�]���*u;B~#��S�>����d=�Waǉ%y�h3��K(Q?���$����^N��[�Ko����>�T��r@�?���8�H� t.K)״��	��ƛ�&�x�[����:�<mS~�i��M���~76U�w�X��q�9��1K��i+�#��,8-�k%����p�iO����d,��KW{�V��q��j��̉O��}�\���ou]�%w5^Zuh����*)������Ti�ή0��Q���H7+����Ȣ�|i��^v"5ȿ��#�(-Jf�he�_��J�e��r�����
�,�醵6�l��5bE�І�$8���n����rD���&�X��'�m����"�]� 2R�v�l�H�	'/I��~��u�}ic�(�\E5�u����!���09Q�OtS��y�@4:���!X"��O���r���B�{ö\�t�oK�!k�w���i�V� ~�*tM:��[�O%�
+�����!��X>Ɔ�����$đ�I�q�+f�$��/��ȳ?�oAt�Q7��d��gE>ͺ�/\Ј�m}��'�6�c�>ڗ/T)��y�1�ۯ��B~qŽYWQ6���!�a��)�cOt_܇K=]|L�����o����6��g_<��Jq�����ގPn��C���������W�N$��p������Cz�24Q�2�5������>(��ˁ�e9�J�@%׾'\ΰθx�'���(�@1C�ʏ?S�
�q�x�2�d��A��cNJ���]x�	zr���=�"�8p�����s�X����h���<����n�J}�|7J~Uby��t��Ps��p���H$Sq�S��N���M�Ż?	`n/���r�Mi/��-[��{�"#�_��Cz��՚�O20򌤬�y�s5���V3�'���+�@3*�r����������O#�pf�t`MK��#��3���/�z|ۓc�Y�6D�'�6 �聲�>4-��+���	&%nl`���[pA	�IݶE��-�f����w�J���	��t���Uߋi�:�fR.-����u :0�h�x7�1��)-�s��j�@�K=�=4� 
�=ӳ�u`o|�V2���n`�����3��,'7y�,|b+�}6=7{�SH�s�PX]S�.�x�ac�0ߐ/����3�:�Z���>ZJ ��@�X�ўbF�d��5��A�*��|���T?�����>E��P���10 tw��:(3��KB��'��	]��Y�Ƭd���Z��N�ZB�6���,5�]�r�v�{�i6����b��%�=jƊN��z5��>!�#��*J��Gl]�|��/Xc){�G�I�Zj��f9D��ڍs%ޛPIo1�w���wM/��t�9����q���"�">���O�� �$�a>�� \�9�p`��E4f��p!e�a��w>O ���A�,���\]"��z����m�#�i��J�6��M�;7�:�ʐo�� cXJ����D�t�������@\��� �{d���P3D���I��3:%jw!=r�'��/��~�.���\����6����0{�30����񪗳�"NPDL{��\�����~�q�1%�ɿJ{ ߌ�s1����C��ͺQ��I]G���� �ՎN`"z��h��V�Hb�������
��{I�R|� �W�oѺ:�3�����(�D���h6z�G"��*�H</�M�����{-k�/����㍸��EɃ|V��2��ף$:��㬄�����Ô{��$��v�#"&k�|j��ހ��#��Yr���y0���Ag��U��!�l��8�ݰ�G�J��̢���ZR���[��n��Шm�@h�g��
�
b��3�������ơ�K-A���_��/������&-���=��8�غ��Γ�{�c��q��u���.{ܻ%q1"�B(l�t~�O��&�w(7�d�ƯY�ؙ�?@J�����X��#�i�ڣ yL�<P����VJ��EzO����-"�l�b�&0T�ۦ8;#�Oe����in�s��ϱ{sE�y+X=��f�����)_�k%���Ή⊯�T��_tg���h����4�1瓟$դV�xȜݿa>Y�X+�kc�����t- �PZ�| �7C�ēL�v�؛�z$nx=��_o��"Q��f8q�vث\���m�0�}
g��L�D��t�����X��;��G��0<	S�y7�a�^P8rw��1d%
(_`�<E'��z)͟�BL�Og�8�-#Iڭ/g�YiLB��D�K�t�v1� ����5��؃��[ү;���m�1����_p��诗^|��L�5F].X	Kq��`��o5�sp㸂��Z�1~JȀ�e�P�=�C�]��j����Ե713r��ו|����%|��b�9������O�y��,���w����9���U�a?'�ۍ��-��T��H��H��D�N��(����_�v���!4 |H²��*�\L���S�Q�`/�m��Ƃ����2���
Q9k�I�m\{v���d�x�F���c�������y+#�";ث{���7av�yO�2� ���N��t��lJ	2������`�@�O �ka0qz�ᄃ�8�� ���`b�ak����P8��WiyW%�k����K<]�x�I�_���X��;>)Wמre����%��S��H�y�r�̇��c�U�T=w�/�E˝��u`Nj=EvbLg�lB
��UF?y������� fU�x/R6md�\s��m��dcC�@�89\$3O=���۟@6��)���g���<�T����q+/���|η�y��|_��K�Pm�&<?X��q+���&e5"�f�癡A#��@�����4�%��ֽ�����n�"k������@8\@����"V9�g7��f3u|�C�Lǅ���M�	���DG�ʑ'��q@��KC��ȡ����m�.Ϋ��6�%}Fث�[o��d|,4�J��O�$e8w�=C�=@�7Q�nP4f����9��IU�8��(WH����R��!��.`+����� �嬞'��&̊�'M:�"�<�/fE�Q�o� �#7���0�1�!LU�y���>:�q�S���b�ny��gW;}���R��c3	3�C�N`&��ꛯ�� a�>��'8RSS�KI.�e<wtq���=�����^�kq�l4UXqa�;ȂT{�����
[�>����^v*��0�o�4�� C񬌎�������@ǈt�2;']2*�k�9M=/����-��@*Y�2�#����YkӮů.�B���_��$��3���|�6�����7H�ė4G���ѡn�JG�[��@d��z�X'������A�!��u�:����^�}Gx�U�7������H�R3�QH�"�߫q�o�Ov�t\0��TAG�q�-�c3)��}X�F�k���8$��Hɬ����lz&p3K	:V\y��}�;4�">#�J�"4x�*p�Yح�p#�LH�i�w�1QH�=PyQ�L�_"�*_����%���w���뇋Ra� �9��\u?L�U�3�(�
ٸ��y̗;�N��&���B�H�i�6+�BvJ���"�������y���:��XT�����u���5͋�o�u~%\�(��(:'6�j�O�A�i&&+ǅ��/X�����
�;/'!��E?���Lr�P	��3O/((敌��W+5j�x�3b�؎0�ݒ��������aE,���ͥ�C*?g��^�(���Iz��翙�aSkפZ.��>Ek��q�Z�3l���rH��|'�3�%7�{���p��k[�q�q��8E6���Cyx�O&Ȱ�H�a���� ���N�`�;"^�\j����)��c6Ԋ
�ta�=CSK�S��AI�D�]�c��G���Ј���<��5b��7nr3%�{y���N�$z�w�$�׷'O�,Gn7 ����N���B�p�dȟ��������r.-�-��i$�{s�Y@+K��T�d��Zds�ar�^��n����?����@��l�
1�>g~��_�����q��#�y�Ɗ{b[����'���t3ۈ�K�|��b�vL�7��Q�����+S���k��i'�W���+���֓�U���xc3H �<��o*�����5ߌ��Yp��H��11r��-�侔�2V��fu3���!�yA?15�[a�R��Q�
�3����K�<�:�p!Se�~6p��r���b��C�[,����ݡ }��7!W�������iS]�T9��������������~!�˗��y P��G��`���[��5�4Z,w�y#w9kS���0+W��oO��1E P7��ҟ4{i�;�rB p�&��0b���9y��>Mo����;B2�g��9�����q̓�j?�h�̗�4qmF^6��|)��2��z���y�*F�G#��s�L6����J���>��O�gL�}����H��j���gu��Du�7�{��D��u������F�*��Ĥ�^�w���}�ɇ�}��F�f��ۊz�[p��Æ�r�n�H
|�����c����*jN�q���@�{�%P;\���"e���:��#�͸Y����)mM�8�l���2�`���)&���0����JP�NO�ҩf� '��RI�=^ۿ�?8�P:7iȴ5ST-�Y�>�ae,��d����I9������k�$�b��?W�#86��j���"R{�4aΖ����J��V��Y'b	�!�\������1S���dĔX���cs�?vة`~`�E����⏿�f����-�ld(�#�Rh(��j�~mWr���kV��	Ӥ���3�]��F����	��c��	�v�^���ȟ��A��f>�i]p������0�C�e\�o&���V�x�Β�%^e��Iڅ�hn�=`����͂[J�ӟ��9t�iI3�;&7,\O�����r�e���0����U��� �k$v��Q���
�HLI�c����'�1b2�ț-�*�����9�]�C;u�fB��F��n/�e�O%=j`P�"EQK��f"7H���N��)�`��u���$�p<M��q��%��T��$��M�ߊ�x`�xM��c�ZqԌ$�/�<g^]���e�#�1�DA?'^�̰�h'-���v�/����Ӏ԰�3s�z���Z���r��T��#wI�*�~��aSN�������2���q�,��@h<��PW�@��6��*��I�pr�%y .��Ch�I�G�]�I��Q�.O)z���Y�G]�����h�11����õ����w�bA��n��a�8�T>Lݍ�-V;F`Y�ѝ�["��X\*�	�YN�.��~�α/Zcd�����&���_�i��9�l=��xR�د-=&�7��="T⍮�q�M斎�&.��`�tW!��LL�_�Y����k -���D&���n{YRH��,�?i� 6El�q�9��������Mϳ�O��aN[ˆv)�#��~P���p7;����,5�>���^j��/r�% ��@'-��\����#�N�(��Ҁ�*P�`�u�ckїnL��>��k�_�S�W��;��7a� �:Md%6��hI*��'4x]�똅���T�zB*���L�<!:vl�R�DRd�!.Z��I�%�"�NSJ�|�a)`�Y��6����oz��׎yhg_G��v	wi8<��Vސ�tӴ�4��Wd(v�a�K�l��@���\R�T�j�T����s%%��rA߇(��;�G[�:���~�w.������rP  �
�}��c��}��S�f���y�q�>���aF9J؃Xz�S�MD��Wg���jM�`�l���8QI�j�$�2���S��Z�3
��wl��N
\����rz�
>@�L�JPf���7�t�VFiԾ���A�����K�Նi�z!b�f
o�a��}-�	2+a
,�9���?���6*��M��v����nʺU7�-Q'�ǥ&ǦmH��et�����s�:��/B�kB&��8��ǀ�ݺ�G
���h�ll�=~e.������#�:L[�	�8im[a�Hϔ�#�-@:I��]�5*ĵx��Ը��\��mciD�`�z�ݻڱ�REZ�+�2}��c�Ĉq`�؈����q�B��38�b,��*�*y���W�u��js�Ő��׬�U��ЏA5�2)��0�KB�\!���u%� �m\�6�����N�ܰ�ϚA�2��q�yHx��x��%REN*�!�}�*L#%�����M����̿�7yB�0�ۢ9���p:�C�!�u�[]�4�z���b^H�P�=���m�ā'MŲJ(�jV�W�C�~�ۧy&��zғ�O�F���b]s���&�
�M��P�8���Oa�;AI���_WL�>�L��u�ǞA4YU�cT7� �(�Q�3�����'��f�Z�B���0��%|+�4j鎵�w��l�v��v0���"ٯ%Ҿ�e��,4�+�zi����&�>.�1;��
�w��2����gFe1R0E}�a���̭��w�ķ�X�+��O/���9�Zґ`f�2�=�����X�璼���y���ŠRf�>u��:����_�	L�V*Uth�g��������.0 �p��<�>�!���S��N��u�9���Ý�LŪ��v%�K����R������Y�mĜY8�ٰ�vũ�@���)��@A����YLR����Ӡb|o�#�ƱUs��q6f�����ٵ�E��%6�rh͠*8ˣ{0�_�b��f�b�yه߁V��
ц�.C��K.P�]3H$���y�ħZ�	�=Q19U����F��������ɮ��Nh0���R'�Ьql�]��e�q�(�}T���u@���*�g����{)p�`E�x
�8�(���_�RղHA5�x[���߸Y��Q�88�Eħ�!e5�����0����aj���5S5?��A'hÓ���Kz�g�%|*cg�l�؃��k�+�L�\�fK���P����#7)�1����p7�꼵ɰ�T〤����eɩ��%l�'y�e���,.J�X�!yʽz,��X:��~Y�@�qß�H���G&���������b�����z�l@���m�q�25[&Y��'WRg���l��K��hB/d��k[���Šz̩[Rk�B��y�+��)��F(��hI?3-R,�	�WU��������j
)��(�A�
��E㿏j���X��&�Ă�h1\�{,]I�UW��w˴����7ÐYz$���'o�ƋӺ��rE��]����$���p�G.a��F1n&X��lc�oq|�{��J42�*���P�Ke��$�[+�P�5���Cy
�;�
pu���#�~��:�4���Paj�"Ŕ4ށ�9��ِ �B��U�j���\s����Vd
$ͪ[�Un���/=6uW��]@O���y8�ڊ�EW�o9)�V���t^��]j����ˎ�7Y�who��d讶�%-���ds�^�R��+��נ�k����GM���(�Y��\#���ΝAǎ��#�tF��B|���![�e�!��\��F

�j�Cy6���hV�I&�:6Hؽ��w�`��hg���FIӍ�NЬĭE��K`����M�u�5��؛s�U �2?�2a�������Cw��\|;��ϛ������6�hE
>�J0%r��@uC�J6�m{��3#���=�?
�&��σa�7x����k�ǖ��ì�@:�`�"Kf,|�ʇ΍�����8�qZ���3g��8���K�P�}k�J���)�������.锽89����^=��p<�W�
)�1��xj\Ǵ2���4ޅWK�a|&;��̓�K��ۓNep���{^h�ᔢ��y�86�'��K��߇M���r�8Vև+��듊��}�A�dq�ꉔ�~]=.-�\T �g��X���D�����V)I�x�I�U��r��τ���̈��V�򂎯��;�f!��ӗ���q��e��1����ɢ���3��}��j6)��̀��B;"�d䉄�5��z�B)�o��K���ۼԕy.�}ܕ�6�e��G�a�>йir�i�!m52����{㲡`�p)��\$sx�WT'c�zGKn��J����f��v���JO#z�Ul[���a. �A�������$FhO`�v$r�9�n����e�Y��r$�Cީ�^薖껼B���������]�?;%�W��Q�����
3T����;��ʓο�/�.�u�w0a�қ�m����Zk�����q�|:Í�J����BdؒR�w��:SvG�.�4��|6��DvҞ�g���(W"o@>��Hɂ670?6t�RN_,6ߓn�K�E^�$[�`�0�
�g��htF\�(+Ƈ|�{�7��Ow&"���/=^rW����RŶ�ch}uQ��FN�cf�2��GPxӾ�SUs��%Y`�Ro�@�]Ep:\m�Ԫ޺����U��l�[�6�L��qY��3w�(!Tԙ<M?\�f��F\�pQ�@9m�%왅��Ħ�v"$Sv�6�?E�Us�+�7��fu��%�4��*@_Q�H:�u�J�V����󶡭U%Vf�k�&�����7<N�Ck���R>֛ڽ��]�f��
������-��Q�a��fp���R�x��: F4K��^І�M	D")d��6��P��{�¨R�s1�	p���ZV�p��Tw�ۆE���W�Ul�M�V���.�B����&\�M�L�dl������~���
�/�+V*�xqԴ뚄�G& �iS.i�{�Bf���m�+����:u^ 7s�������\�r�"���;��Y�5�^@���JH����7t�܎h�C����I��{�bA���}*�pXQ�z��ϐ��sN����AdHg��B��hk8`}�"(��7.;���O�sK�l����s��
��k5��-Ӻ� <8�z47g�5�&�����ڡ�
�|����+t!(%�n��?�1��y��N�R��o��{�m�IGO-n�G��Z#`�یh'y��P`�zj���͐Ã2SdYܠ=�߂���IQ6'��򰧁j@
��]�o��K7�}g[�eH���N��^7��`��&E��ް�)��o������2�@Z����S�E������R�0��n�v�N�2�	�wA��}�����%��y�
�I��]N[H���:´�1�������1L�b�,�W��۝ر�"�:x�����ʼPiO��.�)m��������b�<�f���/¿��i�!a��^��PT.���f�$;����z7<l��K�.���Bi�F��O(�|��&��R��7���H���>)xfy�T�V�R���v�W��=VI��`=�<&i4wo�}#������'��cDUn�3�Q���@g���g[M՞;���:�I=Q����!,u<�R���eN�Q �?0��T�J!�>sZ�7�	�����'�͊�J��0���y̩�C��9�<�b���g��S���vo �����yR����P0s�[�N�S�"�H�k�q��$�p�D�%�92�8�oBYU���~�
�Jh�=y��Í�ʓ�$PD��G"@�g�W�y�ާb��Z��1捋����FH5?Tw�,���3JY�<]��F�;�=)ؿ����ak�f����p�~�s��-B� @���_	�|r~��!ދ9\+)�(%ݔ�p��7��j$U�U���"���B�g~��e�9
��ޓ����.!yL/K���>��;S����p=焵�1̫?�c�
��En�����h|7L��H��II�ur�[���&����M��n4�����[��v��b1A ��?&)p���u��N8,,Y�r�S�e.^B�9��J,��g�wpR>�}��E�Ī�P}�:��+?j��QK��fJ#�{�}�Z�&6{g;���U�J⟆�ϦȨ>���/��6kv3�Zhyc*�#Ui���sC�:a
�u��T}o���},m�YX�,�
U^���y�<ݤP����)��2i�}�ęF�`�~�O�^����F]g$�&����[��q+E�o<Ջ����̢A{B'��k��9]�����8�>�o:�&up�b#�!~W���S�Ֆ�<W���Dh�Лzf�㒷;kY9_��~��ة�5X�Uz2n`�0��%���Qd��r�� ���� b���F��8�ل'�Tu�����(۾�1��U�RW��qL2G�v���
�,��.��c�C��f�I�vZ�c�+���Ƿ�H�f�a|�c~ǚ���ڭǼڢ�~�\�`ٲ+�ڶ��hm��=��[��vP��Qa���}G!���$�78%C�׍Υo[�
/�Y���͟��H����P���XۼL{uZ����!&����^kֺ��TX
���@��O����^�
!骁W�A��X���i�;A!O5�|����,}M'�Q-_�7�R8C�ۅ1�;��Ѧ�i�]T��[�\�08/�I�)L����q�O�aH�; ܥ�b'�qL�F���]��ߨ�+K�sU���JȜa~�Lio�k�^,C�~���I���4MQ�̞	���7
j[�hv̵9��}��g�'G�����
� ���'Ty��T���w�e:��Qm�w� �O��2�&�U�XQ�G��NM�'��SK�_%[^����tZ�dx����Z��s{�[���8��sz�:H�ď��"�8�^���6}�T��b�}��Ɯ��Z}�U@v�`&S��]Y���Г͸>�2�泤�M�6c��ќK�����^�":��:��<#��P�+����lɰ���^������s��_!����FD�W�~y��<(r�o��<��%���/GL�j:$�*H�ꤹH�	�pQ�7�؊�]�tB>~'�����d,UY���҉J�;Z��Dr_+-9g�������+��x��Jr�&?�(�ꚺ��F7��»`��}Ѥ��%:_>W �p �)��e�g���xP��)+;�W�Z��|o������b%p�b���s���U�C��)�����;#¾���q�#���VN\!��S=(@F�lٸ��ܟ�X�v�Â���*u0����t��Δ5�8W{����`��;|v�A?��w7r��p�,���o-�y�����'OsM6694��g`�?x�p5B���ӥxƶ��V��'�|g�?�L(��,��I&����9ȋt&����>�'B5,����KF�	��E_tc��R�)M�ŧL}���P�����J�h�=6Kt���I��H~�sГN-篋�;5��H��P�Ty��w��b���x�Iz�Ĺڎ�����e���+���7�VA��0�J�*D-��B������3��q�:S��p�>�:g�?uM�3-$@0�Ӭ���2�7� �=�JX.w*�o��+d��>����fp�m����أ�#ևpcR���LVӬM�R�ػp�`�)�X��#�|*� ܿ����ѷ[�� �<|�`y���"�����+���v �s�*8����ebi���~^�:�7�<�@�m���^5�p:DY�I�:?���ڋ$`�k��s�@����*�×4q<���/ g�T��qF+!��@o8�c��z�ĨO������=K8g�c��͏����ͮ�능F=-W��F��`[�G�7���K�oz9��»T�?TЪh(���f������"��=��CwK�����Daz�7�p/YV�!&�dU�c���i�@Ԇ��j�D}+x���N��`J2r��� 8B��t�Q�I�'~�g�'�E�7X�rғ���/�b"� �b�����8X��j�ku>b��bK����r�d�ڦ�+��[������$�xp�C5�%��J �ޞ�Y�=X2쉴� ;���M���C�(�L��:��"���Дwy�L5�7�٠�1���l���l�N�"���w��=�]�r����W�NFP��d��Ŧ-u��s�0��.��K�DfU��f���j���vcw�$������')\���c�����T��`�>hI̐�ɺ��"j�b��m����N-*��L��L΄U9�2�7�
H�[�RU[6�:2C��zG�_��O�L�H�8�N��)�ή҇�'��L��K���!W�8���j��ON�9��#��TP��ҩ���n�oշ��uV�_��vm�=��;6A�'{�:vl�P�B�B���ƅ�jZ�Z��Yx�g��.`�b�������޴;�54��-�Dx��e�rI("��OJNa3VZjb����k�q"<��\��-�r��F�����v҅@d�B-��l�\��|�0$+�G���A��	�=y����_�T�@ž�@`�{8��Y��-<?F��J�r%������tqo9��y�O�5-�}8�6"�@�r}x
���	w��2��V��Bm�`��έ,����%�h�X��Ϟk��h9�HA�� �SXq�,|@!H��F� ���>�3�ǩ���h�lф�Z�jg~���I��Q��5PY��	��^�5ʼQ�%����R϶�6�����a8i��D4�����I�}Ed��A!�m�4@�"ԝ �ZQ�@��a#W[�DF�F�y���f���F��UJV�iL�P���np������/������/��9!���r�9�S�xd��|�g�m�)�\��9���!%�8���<��x�Pu�p9�N206�},>����{��j�x��n8�ʩ��B��O�mq=�yC��&b�m
s}����g_�iK\�1�d��S#a�dP,�/G+�\�R�F3ew;��j?�۝�ܿ�q��/�Wu���?*�F쳏�q��pg�KCa?v���o��2�3-�3��]��]F*��3,������Xď���Єu�mJ�%U�y�\�#)�q�EW���E�_��)@�tm�b����?��I$��0;4�u��8#���8�����#��ϊ�5������/V�P�q#�R4�<q㪺ؕ U�Z^l 1����t�6?L��އ�A�Hb$�j�� r\H�U4�i>���9PXp)7Ƹ@�ؘ%>_kzDׇ����㓂�ڐ1¦�Vb]O���g!⫽�A�˒H���	��Z�<�N)�|��i��V���Fj`��`�����D~�
��U�	%�^�Z7�O$�B5��,���ߨ��,o��Ly�s>�c�D����<�:/�n+(�88�a�Kb#�2��jE��J�_"J��`���a��V��g�A��H��7 �Ckb��D�FM�kٯ��\T\V�4HRЯ�c�wGQ%	~�r���z��%my��~�t�M�'�r�k�a �U�t��T|ɋ*��"�X�>��\eޚ���F��~��8�����x5��4��%�Ľ'�xl(vI���n`0	$�IR��^c͟��KNRE�[��U����>��Q���Oc�n��4�M��[�왙���B�4i��Q`�c�^f��]T����r
��Ƃ�ܴF�Ɇ������+�'d��n�:�4,�s����͹]|UPZ�@h�i�^��T�����c�?#m���d���z���~�JLB�R3m�T�A�^��T�R��n��^�|�Q�
;7�p�n_W-�8�AVNM6�Z�)���T"����Q�vh��1��r@��y�G*������}#2���P5�u����q��c�(���Rj�F<]�2ED�;9�[j3B l��|P4�?����Ԇ��~}<@���n~CS�ח;	4YI�ٻv��u������',�~孻����sإ��:�K��h��������bz�������К��m��(w�:��Ί��5�y�X'���m#���/�/\˗��S$m=�8�IGeȌ���ѷ����ڃ{h�q�!�Үe�Oր5��s-�pS�M����_[���Y�$e�{�":@��0O�߷� ��)��'��6ܚM���jjI��=b��٫�R�؆Vm|��F��W(9 �k6\�*�����	�W�;p��ȋ��z��V��{g���ݬ�Z͹G��l�ם���f����%<5�|�O�c�}��b֟�V���w��?��Z�\e2��oڴ<��m�_4^��؄��p�cq��<�r�C7kY��!5���ׂiyrg*NK�y؜p-��Tb+۶�|d�tq�*���2�;=#�He1o\�7�I���r3r���vU�<0:~k�l�0��!W���n�GJ15��*A۹�ǖk����"~�����P��[�)��,*���b��X�.4*;)F���s=����ğD���z�_�ͅ0R�a]���{�� � ���U��͏Q�Jp,^T�ҙ����W�k~Һ������� ���~����1��`�"c�}�~$i	�\4��⃾ɻ���k�e*�b�.U�^�A�ۅ š6�m3��KT3�cw�GQ��ne�����\ӎ>�z�k��JW�x��wݝ��U��Z�5�&E}���B�6{�O�H�������%��wLG	Tf�*�b9��̡��s�;��E�0qb�B����Vg�;�`o_O���{lɢ�A%_��S;wݗ�܃�/8v���!��*��(���3�'y�|ʣ�Z�6S�t��>t�W7G���DGC���sk[��uI��yF�0��3�3�'��2�Xl�6��F4F}��jA��Ad#2��%���oh#@��h��p��ebP�y�d���c����)d O$GKP�E.��Vճ�Wb�޸�V`x�u��7���:�ϙ�!}J'@�Eȵ$��f�%k�X�(�?���JN	�+��ͼT��#�D����)f�����2�X�(�鬖pkk�\��"�d�K����{��|����!���-��\ԥ�|mH�-�"��-*j9�>th�Q �_��m��Fxz����Ú�@�I���]~�� ���J�m �.Dh��NgJN+�}�I���T�簋�_��N��O�x�g5��j@��S�ќDyy���7O�K��e�$=�^4b?v�t��$�2����b Zⵝ/��5Hp48�a����K�B�^?�>������
YI!�r��Ԡ���I�To �Sr�K�{Wh���7×���.�蔲�޸ �H��Ӽ����|�ڑ�Jbh�E�������XTpױ:4��CF����e{ d�٪��&�S����6r�?�*'��~;�5�W!���.�.D�.8�ߡm�6:E����v��D�#�G��RN��yv�go���1g��ű2>�͏�U�¹b�!�j�[gi��=�^v����Jnk���q5Z�q���u�h qP'(�����e9�ܢ�)"Z��)�%Y|xL�� 9`�O��3;���!K�3zЍ�4��Z�s}!����&�b7�A�
�ǝf�?�O���b:�S�%oM��_�^��#~q��e�L޴����Z<�B�Z�P� �%�`�1>W�D�嚕
.}�ѿܤ���}
���I����7&��*�\���Y��B�?6O���=,d�0f!�\f���2�j�F��� �l�����q�;}v9��tί�3��ˎi�圬&b��E�Se$�]W�=º�C�b_��z�����}|a&��a�P�	�$ax[۷�����R@�lvP�A/�QG�6��	�֔ {���U>�IF��4�k�2���ܱ	G�a�Q�a��l����� �(��|��!7RbG~��� N+ҳ�fQ��(|B������:(2��L�I|\.8DfVU�����_��po�-��j+ 6cn˾��ʩ��6o7-[�Rf+Nװ�BOT��,
��0�	'.%+b���AT;��A09I�q���R����S�M����;rۅH��,V�|-��-�k��	�{n:5��~\��f��N������j����5=�W���!�<�0o�;��}�|��^>H�ܠ-�SC)پ�&s~U@:>`�~�d*9s��d���RԻ'{���i�_�A{�=����[�]�8#5HLVq�-��cLV�7K���XQ�A�1�پM��"�n�^5�B�w}��V[�����]JPF�v���<��_bV�OCq�j"��*�jڹ��c8�m|Шǂ()>���yq���q;�;?ܞ+<Oj{���I�J�%�r� y��.�Њ���A6��K��W������e�A�w'��O�=g��}k�Ozb2ug�.�X����Kx�M8Z0�B���x�۵l�����E�~�~.� ��D������N
f�#�Uʇ���/t]�l6ʬ��S��<����$�O�@y�3��C$���IU���0�hn����Ze'.�����b�&E�B���2�x
9��QkO`;�dS�э�����\+Ʊ��cUj� ����%rA����x���o7ژ������6��|}S�Y���I���s�p���yd�|C�-+�{��>^�����g��˜�4&I
���J<�\T�R0fUq��Ä�}yQvJ#�k�Q�q�s/�ل�u��54KL8aGҊ��d�5���
C͐K(AA�(�%�
" Hj{A)X��4;"|�V\�̈́��-{�m���=��ǂ���(�O��E``���e���yG�&)R/��'IPd��ֵ�����(�����h'
�� )��s��������5%m ��{�,�:y�{��U-b�k[��SI��{��d6�M5"�1�\���My��{z&��	����IjF��g���۹p���N�E�PwuI�,�<�	'��uEf"Ϙ�f�'1���~B[�7P�~���η68�Z�vsb���}�l�K� �B�-��]R�ơ4����F;�WX��]�Mc-ٷo?�������m6LC�m_Be��-��ʍ�"���t<�%P��L�.`��#~��_GE��2/A{1���nT�����l����ۑZ�K��)�=p�]D��-����� p�� ^�=áz>��C���ƴ��$c'�� VC>H�a�6�a�:��X.��(^�[�H����o_������Q1-A��ڦ�l٦o|��inc�gY��gF2;�_�w�/ϓ8H��f]��F�Պs��'��-�,�0�����sr�F8�Պ%Ue����0��Q$����*���o#
��L>T,N?�]{:�[�\���%��u�R���o�j��<�W�����n���`���r|�|)�m�E���R.��& �wl"��aS��C��,b��Rڨ��y%�:wl�M(?jE`�u[�>�Y�+��j}	�Jd�CV���nẏwl��y�7�c�;T�E͊(����sg8g��vtV߀Ѡ�bii�M�6_fXo[���|��´�U����[j{��Z�eOh"A��q�)�w�yMoNJ�\/L�zVT�J�-n�i��E?G��k��k�g6`��!-�f&��iM!�5C���.���J�n�n �37o���̦4�f�a����h�f#�GS/���G����$S0UŒ)�kp�I���[MJ������8�7�x�.U��tP{�)�w��%Qo���`Xe�����c��Y�N�*{�6t��8
�� ��h�Fޮ�yl��>���y��Q�]�"��Z�p6:��O���,�,�P�q��,5D��_/0��J3�uJ)s���&9��K�n�?I��΂�r��,�.3�A��U�WT�P��3���I���H?ͬָ8�DR��Y����x��o��-c���k�Ŷ���vV'`#�x[�����Q�>�k�P�6y� &�v7���+�'Y�m����eB����堑������a"���L.Ё
J엱KSa�!��됈~t�e�u�I"F�j�+6Qt\�c�vh�=�]����G@\*X����Ou���b��NN3���xbꖏ贴Z��� �4�?��)��O,D���Ց+��/US>U��ċj�b-v�dE�����3���O@`�%�� ���h�vN�u�_������?��y�Kz�/�sƨ�#�4h��-޸��CC�0����l>�$��������,eh��0u���S�1.U�(�[3fX

p�+�ũ]��@�HM�`Dt�ICs`Ok`�x��0��0�9O�a�'�[	��A����)�FI?��E���V�$^U�|��M���15:D1X����&q`�ll��s������x	$�p�[Z��E�r��^%�mq�JG(��ah��+_{`�m�vS����9W�HS�Y)z_�,|H������XJ�.~���?ʀ	�jQv�_)f)w��#��:�����Qx��1V]k�%[�oD�M�KWHT��to�4�(K\n^ua�W��4ݚ��~�ٞS�q�S�cw���+}�y���E���W~��X1��
-<�U��,�=��鋾z�eV����i��� m���o�M���M6($Y�~ٮE�F!f��m���u�$�3�rL��z��>mC]��2y��Ȱ��Z#�bn������W��҆�q8�{.$����~6��4��\^�AyH�7s���C��C��)P�N���nx�[�7ʹ��nNVi�_�����GP:p�\�m.	��;a�`���_N���[�֭�u���l� �ky�?
�P��f��Y��6�F�h��	��TW�M�G�C2���,_z���)$O��[(�뎽U��c67:�C$��`:��k��٤}�_tYIa[����x�=�TS?��h��Q,�=���J����D�	[�H�|j��v�1�p��D�4��$�G�)��o�S�G�G#p��H��3�܍$)�9bH��񷾢~�g�0+��H���ye�N��<YX�ɂ��T7��Y ��"�~^eU q�kڙl]���|D����U=��kR֮V�+�u[]��@+c8$=�i��Uм��SAz�}����E5u��~"�V<��c�&��Wl}�U���?�1"����%I�g�{1��b�&�
|�oE��G-�f��~�AV�aaKZ�:2;MY(�,�k%D��08�'�
]�o�Xߜ�<G���oX�TJ���к�m_ p��l��V����:m�!��g�5m�� �An��&)�?��"��Y��R% |�[MJ����Dd��m�!�#���H5�p�?���B=������0Q��S>~���	~DSl����n��n�S#� ��DCf�7�e����B�VJ��`�p��2�~��\����bM�A�����b��G���9m�L��W��# ˌ����L߬��;�o ��"w��j�9�P�؁��e$K�ɜ˦����J�fb#q-��k�2&��̻r�;���ur`����t8T�@��y�i�*k�{�l	����~yC��j�<:&�_`��q̯�n���ݚ��$�o�$�5�I�+q��2�=N��l1u����5�v�^�C����*�b�/~��X��~���X ���\>�)�n�R�yJ�aeML;*W�g�CH'����d����G��	��×)�$e;dZ	�{;�<YBT�	�j�����[9HqE�C���9���P�T@�X�9~�_Aq>��/3ɉ˴e�|'�O�\p�-DcQ����4�*�u�ɘs2G�i/pJﴯ�/�p6$rŤa�o�/�Vl����|�/(V�<:^���LVg@����.F*��+y�ef~5D��#��ƿ���	��Q���פ�}���i����^*���q��"�Q��O)���3)�n�P�0z
�7S������η�ZRLv6S3 ē�#���bp���vا.����G� �D��S�@3B\�]���%���? ۏh-�t%J͡2�p f��M6`:.���7��n�z,�,=��琙������<P#��.r�A[����l�!�1��1ׯך�v�K��<1\���C�:�g����qg��ݸA�� ��*sph��*�H��.֍��h��<���|�?d_+DZ�V�Ӷ�x񭴈ƹ���\�P���*M�X�s������~\�'4��#VF�n��x�=�Bґq���z:[��m�&<�mjs|0�!cr�t:�v��SR�Q��坕�����@+g�}�W����� י�N�z=a5�s������ gCsUv����!�|�����1>GC'�
	��}��'�,P����X{F� �P����r�f�*H!q錕*�J��k��7�ay��n��g�eS�t�OMgyH�,�xHjT������q>h_�G��޿�����V�����I�PA��mO�hD������2�,uz�`1+`��	Uy=AB$�y� F�m������_�OP_��Y�Kx0Ţk�v٢)(gb�����4g��cJuFt�;�zH\�ƾ<�JlM5��ݻz&|��u����Xa�z���F�QMm�A�H�'�ƼXu=se�?��N��ר#�4��v�v�n��\U�����q��Q��c���'\���A��F4 1� �^���C�m��K	7P�q-��i�-0_��&�|�+���7�1T�J�R��?�8Qk4<���.����z�f�L��4�����y���iW���v����
������[���c�-��"���+P|��
!��� ƚ4�ϝBߥ.M��&��p,[a�D�?���"��<ͻ����n?	�~�m���&����Y��U�uX�b3�hYı��>�:�@��Al���TҤ#�������6W�a����M�q�|�<�BF�'M+��CbQ�ʧ���f��C9:Z��d��Okh�ؙ�OdV�	���AE$ ��E���	�����gp�?�W��e\w>��(��yn��0�'��7$d��{I�ݬ�f|{!��[��{6��N�x�4��F�u,��KP̅�w1�n��
7}�-���x��63��&��~xt����%��E4{�Q	-��^�^�V����LVmr�Tl�T:�HQ��t
�B�)����a��j����L�@�����ck���w�Y��b�O�I���E�rUN�r�#�� 
AO���gPx���>�&�.5��[N���o�[�!+��u7Ih(�-r9]W���gO�1��4wIV��ɱ��B�S˕%����SP�iQ/� �"᜞�����c��9�ﯯ�pWn� �׌�-��e��!P-�"��2��j�y����W*¨�"_�i\�㿜����%���"������J>0G6ˮ��ȓ�Q،-�o�mA��u"�� �o W��a "W��y�7FY2?j��a֫��w%��`hI�#|}������Kya?3�D��a�Ķ�V�!�>���{��*��"Qڂ~�B��|(��4�xp�)����*�s���Ә��a�m ��?]�?�ʵ��-~�/~�_�|��$f�*?�B��d+n���t|�+�+�Y��3}�&�<��S��Ɂb��~�J>��B���w�)��]�.�N_eĊ���V�]f�T
�d����\������S!�l����Gl;黩p%(&FS$��RXņg[B������D֧L�HBS7�P]RmT���Ak@�Ha1-�v�W߄����I�L�?���ÞiO��5��1k,�`�I�`�dc��=�	D��[��؇nժ����n����
��du���](�Q7�7��7C����c� `�d0���J�T����QTD�� �ʿ9p�X�,׷�B�w�49J[��d���s�$&{7��P^ : <w�~xwG索��glt~�-�p���;jej��F�V����&z�L�M��s�{p(W5�$-�Ժ�3��޼A�ﶘ�~^�Q����U%?gD������q��p~���d'�E*��v�
:�����EC|V���$��]ݘ%�r��;���s�փ ���܀2� ����@���6]_⍤���4�q����M��Y�s�g��{z7J2�Ȫ�^&1\f,:�� v>X�WF�.svG!&�i��BTwW�Q�&�g?��IF����J�J<�0c�w�g�8r{@v@Gm�uC,(��*'׀`G���u7�sffP�k�}x�zЭ{a+�	r[����胪Pk�<�A�`���_��W�U{��Q�.��vA�Ȇ�uL�A! ;;�klp6��甘F���%L����ޔmrѳ���uD��)	f��6��[�h��1�)V '�	¯�"鳙�g���H��a�
��X��q��S�� ��'�sv��N�􎶴^ޮ683揶��ip�x����_z��Wvح�����~��B,z�3��E�����Kpc7�ݼ� �Z��r����x%WV�7��6�788*�rh�#i J�9/��<��5@�\<m�bO�D��[���FBvڤW1B����Pg{֌�x��myx��]M�ܔ���F�a!V�����}�@��5�b�Bn��܊�j�㎆A������5�4B�6��}��[�#�3�bFuA���1�|���]rl>�P�B�7<��VWڑ/����Kà��?�*�����s���a4Z�D+��B��q�$�`]�LX)�Ė���mv����E+�p)��E$�KJ�O�x�o^�kͩq�9���e־n��ZI_a^���'nC(�w��eဴ�	��|��`��39��,N��2��j�!b_�X1݂��P�E��5z����e���M�>�̼ը�[�`'8�e�������@�sv���N{��s}�T�f+�H��͓t��e�A�Sy�Q�{���%���h��8!\�ӽ�a�\o��z�d�?5�͹}Ϗbd��m�e��oNH�)6
��͈���\3��N��=�e��N8���^T��gez\��en��.�5�������Vߖ�Z�#[��V��*fLa��DJ:����a�.�/}q�� ˧ʛ���J�6�P�s0�k�N��~fY� ˇi X�7���%�. �A���A����V�k���/(�m$͜sV�I��&d���n�Apjy����"�b��o�čȦ35�IIшL�J��/G!˧��3UB���,�ƐUsز��Ο*w�\"��@3�M��,h����{��cG�!�N��������᚟�@�l��(?t�J��fX����$��Vq���ו^Igl�#CD
%~3�
j���sە��
��E�/�����v	��"�y܌5�xR$�B�ݺvdRԥ-w��9	�obU��sA�aPLK�2:?�-��D�m�krhl����*�؃�2ѽBu�ҥ�8}����;�˹���= ��_-��6����N�3wbF�l�J(�9�<t+-�n}m�:�҉�w��w�Ԕ���F+�ŵh��G�z���`R*0,�{,V����������"���Z䠐:@Ѱ�M~}��b�+ g��V'N��רa7����W>D#/�R�@���bb7=�5nH8���ʊKe{g�c���#Z�TV�D� X's6�n�����,�Q��n#8�ey�͹2���eұ�ŎU��+S��^�wr������+��?���'=;S��5l��WvmJ\��B݅�B}~v:"�Ӊ__�kz*�i+�.+�Gd��y3�VBZj�}$\���� �9s��D��ʗO���_�.3�p0��@��V��~՞
Z!��n�īH�����a�o\�|^(R��!K�#���Bϟb�U˩�%y��X�f�ʝ���݊��X7����};���h���_����� M�~#�gRYB���7@r�.L��
�e�pߪ��=CdC�B���� ����G�t�����tVA�V(�m��~m�c�j)>,�C�����ԯ1�:�����<�wG'�H<���+>�х��-mEi�OPGi}�F�-������RyΖ�d�*��~��O8��CL���k�,�U*>��)I�|o8��|��=�<r��kPf����D#�5�7u5,�I���۰�hI�5uC�T��\��,0�G�E�ʅ�{���g��q�?=�pRӇ4V�<�#sy=K1�!�n�L '�8����#+���_|���U v����kV�hiS�A��'�O4��˟fɸ��D.~�c��� �Z�8��g�`򐤢E��� �>�bk81�����p6p�j�C�Wy��PZ��5+�!(�j���TSA�8��)r�rzI
���i�3�+c(�p}��a���]�WI<,H蓼�j��ց�\N���)��28,�#t��a�����:�;�̔`ݦ��8[;5�a4��k$q��V�}�߅���>5���}_:Je�JcG��ѽ(�yg���_&7�c�3`�WF���ԏ6�������z���a	�Q$�Tw4����~����ېB����?�C���
��:!�K�^��E�d{W�n��Z��剽H��?U>�K%�y@_i8a�BXU�)���@�9֠�r���C��o�Z;������	)/�l${1B5���1��8�ziw�8�z���S%������ċ����׷���������K[�AR���#�=����h���F2nh�-R�H�g���^���a�SΙۺs+ܾ��{$̒l��­�D�Z���JO5�.[|CM7\��ټ�a����J5�<Hж5s�1F�꩷)���;?�_��b*���`3`��+՟5ܖ'�	�Q>`��6>�5} �Ї����B5�=��?��~��q�<��٨P�S�hVo)Sd���Y�}Ff����w1<f.}��)�w"'��G\l�0q�4�^�5��_��nk�J�틫���u�[���|8�0��*����`�*��xK��5�fRVu�m}K��:k�rd��3�o�#���&��ΰR�]q���h�eK!��D�&4s�t	�=|�>ݵ�b�������Ő�I�½�h�J亊�n"�6���_��|�03���x�����Qԙj$[�����H��Ю�"BI��e��xs�b+��RS"��,�~]�Nm�6Q\�K.��@�>'n~�i��c���)T�٫�LkP&ݎ�r/���ߖ�c�l�J�=6����o+��k;�m�X�!ݓJ�)�>��ľѩ�������|tv�Ѿ�R��h��dWj"d2����ɗ	������m ��+���^7������(U�#D��"������۲���u�0h%���@��}�A=d�2��4f4C�8���b��'pMWv��S�o�UH�o��ֺQ�t	>%Z�!Hvw7�w/_׸F��P�-߭�{��YQ�T�w��C��4��hQN3������׀�`�	�+�9���6wO6e#.��}�!�����ڛ	���xeƷ&�K%�w���G��2�sr�gL��W���}9�T�9�Ħz��7n�Y|�����X0�SN��g�9���y��H]�统;��E<N��[��@�c��;��������x`.���Ax`=C�y�Z�\�5�n�P�H�:�`��TQ{�s��pwQ�5��K�4�Y���Z2��W���D/�ɺ_F�h���Dl�"���a��d2���FXm;ޕu����|�
��{2���Y�E���P5�T\+��9k9��M�K��{��+�g.��cmW� �F&ׂ*:�Y)��sӃ��U Ig�fȸr�Eݐ���@S���|�$yiK��rȐ�s�V���}�yd/���e?��tހ�t�ܩ3X�#R�ȫ'�/�^���H}&D�?�%���n�/�&����EWPhY6��0��g��s���D�<4�)8��ѵ�{Jd("��)%Qn|։��R�4����Ua�W����ŋ�kM����<�i{�ѯ�\3Q:������k�6��Ȁ���&es �q`�:�漢'C,0�����͓aS9�������N�f�lȳWN�u�NK)wI�hCꯏ��%8fd�oӰ2ʀ*G:����b��xtx/�%������h�j����tO'�ng[3�Q�D�zB"�����E�X+�W�:��a�\���b^\� ���Қ��Kj	��>)ו-�e�fҠ�� ��������*��!��L�Ԫ0e��
��Ͷ]���A������I��à�%/]��=rL��j�<A P�Ù�0�^�:��;�!i�����C�R��:�˥&@��E+��hF������W�Zj�K>(E��HMIR�An�����L���Ñ`���p�$�B��M>�+�s�-�)��{�ۦ	�߀ئ%�~&X���kc.��J��p���̿�L�6Ԯ=��nV@wGXn�� pg��t-F�r*IѴ�oT��,�LG�Γ�os��jazv>߶�v��I��gq@�+�Ê�n	T�	u�ڵ�������7E'^C8��N��t=���=��E�>D��a���Q��ߦ!J��]�����\����M����䉽��GǏ��{+�ק�W���]�'At�Cm�-�
�D�?��o.�L5B�thAJ�nM�2#��;ߠ�����J�xH��RW���؉�N�5����iѧV�b:h�:T,���i�:
����zA���1��Xh���!�5+=�S�Y憬���-;h'�:�i�VN*G+�?I6�j�<���?	�q����z�4Z�SK}�l����2�0�+��b1U�2-�(�ڣ���9:й��m�PϮ��D--�F�&b�=x�}厂��M�y�*K�R`T��J�wK�6�G\��Ep7��d}u�C�v��--�*�>1�5f �	�i�\d~V#�E����+�YI%����B��
]��w�-��8D~�I�6x�l�>�Uv0�17�t���}�&�F�&?oa*m,��'�ǙZX���@)xS�3���|��-�,r���]A��L{�찆��@�{�\��.xr⍌;"�"刣1�]R#e�8�۵�g0w���i��$� *��O�zt�?uaO������N��˷��f+�ߊ~���������Ʃ���ҙ9��99H)HAp�1_Ky��:?OŢ�;TqU�i���⍛&�"���H�R�O&�m�����Ga���Bv0��p8�,s�"�63^y�M�a_���^/{�"_�Ǚ�t;�$b�`y�n5/��*)r�gat�9�1���{ѹ�����-�߽����MU�݈��C�a&]�a�Iw �꾈3�-��X���C�31خ%'�.����C�e����
9�1,�wQ��zj�
(s<Z&������}e�-�ڬ��6����A7�+<����<9��tpý�󸰏`��ߖ�c��_e�J0��D�Ě\��h���1�}�ܰg,$��Ī�	+J2vEM�Ņd@e2r�˂vl��l�U��M�<�x��6���g��mBϹ#2�W���H�|,zcwE	I�+~o���RE4�
T}��K�咤^PP2c�9F��CѰ��^w�/L������jỖ��e��T��[>��6vҦ�=����ׄp��5qTu[�uH{���#V��,ʈ.���3����G[8Pۺ��/�y4���R�Λ�ڽ�y�V��)f��\/ס�H��v���%w��;Z]���s�z,���`l�e�8\a��$T�n����JTd�a�{yfR�K�t�s�N��w3'Şm=�)B�k�6����#��L��}����kb�����D�6�>��U�,��.h��4�˗B��B�٧�c��'�3ڕD��µ��\��}����ڿ]s%&5��L�b�l}�4XH���F�+zǷ�_z�����"���<��(�>�,X�����o<̶=X_�I�q[��]�%��D�DBq�kJ�z�c��æ-��G���,���2W ��}�d��K�p�j�����{Z0'�=��� ��l~8�#Ӕ�����:��?J֧	3Ղ��� �5�����IFB�����JЦ�_�e����_����W��9o����<`��E�M^���=Z�`��ع��� ��i�Ы������SUɝ�'s�����o�0���
�TSA��!;#A�b��5�~j�������W��'�&ʞ�i~bd�O�LG��=��.��ä݂�Y��n����Aٓ!<�DV�Cʣ��֒&$I�5P��d�W˛��	I���̆(oԗ\c��u��h���a��S=u��h�J�yN��-Q�+ڧ�����d��������*5#�~vS'3�����`slST�|_�/ޝD�1H#tև����znU�����b�ND��n(}Y+���݃X4m)'�w��}�
�C�R��91�����<4���НO�ue�;3C7�;l��(5�ep�� #㡖���=�������qȟꖒq�t�#8
���)=Z��9�ܢ�d���Z��v�00<���N�_<�<���	�@@ɦ��;Uh9�7������F=�-��)mQ�:���	dm�w;��ʷ�@?�]�+<^���V�Us{�����1qz�G��5��Mv��A6G?��l��@��N�
S	���Gt�/�Ơ��ay0��b�=��f��a�Љ��ЗKN��MR�����/o��\$U�r�.���6��K����P��⭔Jtn���~��/v�5��"�~K��$�n�m����d�1p���w-����4�Z����N%�C%݂Q��#=�rs�D�o��ͼ��fd�-,�!�8.��
(�[���5%/N2��#t6�������&�	���X$O��A-�_=��
��W�E	�SK�9KR��^��K%����>C��.6t������|T�C�]C2t�_0Pq�V���QF$��6c�#�'[�Nz\�|רv����Q�B�����:��LE�m�:�gT��w+�j���G�TpYOL_����S��X�ӽq�'͉]QB=�/G~�����.�|�k6 �5��)�/1,�%�p JG�@�(�P�]����hN(:*,�ޣ-H��K|����$���%�:2%�Y�<�܃�ʁ�8��^qE�	�K��PYՑ���K�ż��5�è�}STnA�`�R�!�� c*&��S�b���,g�hҒ8��}�`�� 4�aQ��G�-����!8ݺnnB�.�s*Fx��tU:9� .��������񄫜�5OMy]�UQ6R�����w��u҃�Mф�G+��� 2T҂ߘ��ly���?�:O����X�����L>C����ұ��������EV��X�Fmf����v��2�a��%�_lÀU�1
kR�;�DgӉ΂x�Ȗ����7G}ua��Pt�N3^���5�;	ˮ��kV@�II���bkh&�#87ybsk��:���ċ�JN�S���SCn=)����b��j�0ߎ�x��Sr{KsC��$ö\�an�#���P���3m��&�"�e�&|��2e]i�������XB���*��M�To#,]��c`�G�`��y���,f�$�{O����/�oY��W�E�9Ի�l�)����nk�^Zu�eǠ�*�씏��@gW��[���}�D�VB��B4��u���k�4����`�N�{���������j��G��'A���/|�Ȥ ����u�G)P��]�=�K��uZ٣���=���%
c��^�\K�3ͨP���k�Jucd���ƪ$�2!��� ����j����]��\W� ���6Oj�j�
" 1����"�f��N�����(�"rh��GQȔ=5��1�>�+��g0�<j�C���:�$��s=�=:*��`�����������d��"���J��d�.�d*l���ԡ��<!qsM����N�&_:�.�Q����ۂ���5�tV���r�gtB�+�n�]�[\��(KE��
��`%L����,���`۳@�[����+�gٓ��3� �@��&@�qt�J����=KcO�5|N�+�cڈ�'�Haxxݫ����;Oda�R�s���
g�|o���,p��RZ�*�4�-{>!�TBeVcR^d�c�FG N�Kb̚���6;���F�P�la�����ϷU�(���R�A��)C~�&Qf�|mv��1����͗4�7[L��ʓ�ښ��{��:x/M1����gڱq��[05�u�� �L� b�`����������am�N,��(�AT�5Ϫ+Z��E��O�s�e��
o�X�Rbj��p�eD��Fv.*tא���4�!����<T��Q-Ң�S��id�4��ۥ��ޞs�<|�7�>��.7��8����}\
���=�8�:>/�N�3�T�:�U�A��,��ʟT��1���4�����ߵT��4��T��� ���:�SĨnXe4�ӡ���S�<p�=4��D�/��H���I�W0�����GbL���������v�dW
tA/����K��r_F08���5��"񜐘��,qh��RM��)d��w'���k��J�v�m�t�e{��pVAxB�x�@:���Ta8�6�D�P�Ȳ܀6��m�G�3^�F"|�O.?��6���L���z��o�ZӚ���&r���E�O�٦8a��G ��?]�[�D ����/PFdʢOD��	��"�x8�SW+�a��"fs7�g���;��"�c��DB��>�4,ض8[��n�&�A����+��`�5
&�<�ƨCd �Etq���H\ͳr����A�D��#F;S%�}�8�q"��L5����{����;z��8}��c����ԅ텕��
�a	^�,|Ҋ9���~���C�/��CGI�{��<U�!6�IEW.fy��5g�6u�7���NEe� ��8�"�&v{�����D�I����M���>��gR�/�C:������!z���&�k�Q�F=M�>YQ�}Rv��!��������i÷�q����U.-��e�m�A>�կ̓Gq]������}��N������7�(��rB41�@UkY)cG��J�:p�o�,Vu�C}����u!%������lvSL,'Nf�9L���A��`�jL��pb�)	�!d�	���Ed���˛�v��*v�+��B���R�i��f����'�n#1��X�e��e�/%�����4lt�37�q�~yӉL�� ����.H�|I<��t��tgVhҁ\��z����j���*>��`C?��G )6yTl~]�%�F�;�+��8�ᛳ-G��4�3In`\Z$��9��_�2N}�c��wQ{g_"JRN�-8f���!YL��F��G����)VIM5��n(A� U�_��9r����o���2I=m�MҺ�w�}��sp7�1EE���u!_�Q�������_�aͮrʧ�}nKp�g*�
���(�@	΄
�^sO�Od�pҁϓ4y�z��9�>�B������q3���6�Cv��$6)�k� �PuŢ% ���i}�t����p��W���02�4c)1��d�/\X)��ч����L��ȍ�nů(��CP�&T���vMA��	��Z�P.�Y�肫�E��t����I��Ӆc�D��6(���f�@�9hٺ�qh�,�;Q�.#6���gl9c���Yc���C�t�Cj�(�ӂ��.7?GY�L��b!���)��<G��&�z�[?�����Hj�iWh�'��I�jt!϶��y��c`��!��%-�Å�ND�P��EnoT�c��*\�|?�<�k�ݹ��";F�Epk���7�x�K���d[������*}�&��=�7,Ζ��(zF���Y���U�h/B�FΏ0;q�c�9Znkj+Y�Ȝ��:sD�Yn=�ir$4�"*a��V�K�~�W�l,,��^���^H�ʋ���m���)�dςܕ�5ɀ<��ɳ��	�a�-cϕ��C�F?
�Ǡ@*d��s�Y�<W���q8W {��x�̷G�Q���Ф/Ѕ�ٺ|����s	�}�.R��"����bF��˨���7٤Q�0B��(��_�O_����w:�6��؊.��!$a�P�՚q)�,����~����NӀ�p��^0JJ���U�+w�?���D���E|�T���|�]��P=.��j5��k�'xa��3�P�1�%��D�g�\�7�d��)�<��2.<��1��YvR�ۦY|p���>Z��D`w�Ңq��Wl؍L�ό�郲A;�>q����HK1=.��E�f�W�`l��)����jD����2�&3CZ����t�A-�u�>�z�UNV�]�M�'z��a�,�`�w��aV�ę~ьSq�X0)`�_@$b�����U�O��96��k�k�`�Vqg���L�oq�j<o;��uԁ0!	S^���DXp38��9���tʓ����t�ݜ��
��>�+��b��6��H9��Q�СlT��$��'~�Ҁ��Fd���[~�����n]�WP�x$>����BS���Ξ.�s^�M��Q#R��^NO@;K�;D��XTQ}�� d�]�Be�P�F#(�e���Y�NBX���;a�F�3��!�4c;���<7�_NWvقRP��j���H����i��������C�:m�	҆>���$����u�L��ǅ�a���g_*�b�#�>b�h�TX�ѽ��0[eܷ�d8D�'���t�~�ZR(��Z���y���t�[������>n���z,y�L�It�3�`�~�o�8|��,BUr�{U>hy��W�K����T�*4��bG�{S_X!���u��䠽���Nt)�	�@�4��f����mDfy`�N���y�VM�)�P��.�"�k�Ҝ'�2B��~����2% /l���v-����S�ho5hߴ|Ad̎p/^:!��A� �uX�M=�6I=�3
��h��@n�x�~]s��ՁH�7��a@K�S[��!�'t�F�OIv��~�PWr������.-��_hb��&-0vy a���Ӷ�{;N`���5l9�|5f�Vb�i��'�hXT�S�]�!/8E��5jlǪ�Dk��z�gDηlP(�;|v�� ��r�)8_�䜕�ڻc�к�4C��Q
��&:��&�U�<��c�#�<�ζ�U(�^�7��*�GeT�U��|�=��=5�5��k�ȟ�
�m�}�5�����(�a.��S��Gӈ,sF�L���3�N� /M'�S3g�a+V�D��UC�K̂���l����\`s��u�#���{?��O�G�+4��(�,u4��%�C��1�_�m	���ʚ��N�6�G�M�P'�7��%)�D��S���74v?��U��]�]�y��ݚ_]N�"���}�C1�L��x~���7{���5Z �����M�"�~��Pق?@G�Nc''vy��7m4�;�<����M&{2\~�KGX�G���tך���LK�iC��N�d�"���C܁:;�m�Gx�X���� �W���Y��V"�l�;#��,��H�)�|Y�X���ǟu^��{�П읧�Z��X���w��{Xښ�hQ����Ѓ��ۓB��R��Q��u�B�%+�v�ԳᜉV�[M�~�@������#2o��@�B�=���
"N�8zSK#��zud�ʑ<�ҧ�>�3E�_�~t��C���*��|�Tw�_��𚴙�}�U�Z�빁ES/��Q�O�~j���*W��-��׻s{�·�~��!�p��e� G�6>�tV��\c��0)������z��^w")�Ɨ��k�`�\�/�IK�nE��Cj�˸U��������c��L˙8a��M$���Ef�F���#ބBV�� ��[��ґ`��pVIJF� �/'��&�y��c�҈kN{Ep}�YaaR!��dye�X���|�m��&w���!w{�Ũ�W��A�^���Nɇ_� $/=�O0��Ďz���ٻr������(.?�TJ�r]u c�2����
i�k���uNޡHФq_����a</�!�0/A	s�Y�Q�`/��B������w�1�u���`<�[W���T`�$�h���u�L5�uɧ��٫R�+jBP�T���St;R�-�T�b<Q E'�8]���nI$e�6B	�}��񦦗�h
��{�+��cS�ӷ<u���6��ι~�&z�Z;B��?j91�s�,T���UIeT�<���.���V���D~��h�;�&�bo&�i���(�g��Ր�g@*��|�Sٿ�p�摮���m�!/�^P���--�}ڄ�IN��aN���(��F��2A��,�<���I*.Ps���@�Y��D���_�M7��~��n���ۃ(��7=U�C����F��4t�ŀl����K`�]���}����pi�/vC���˥�}P�B$i�[�d��֍l��(kg�b{B~��ֽ�;�" ��MARr����E�i�ge��X(ӐK�g"oI���AG�ݸ����Ĥ����#���|�^��A���Ξ��zΨ��<5v�Sq�>%�%�R����#�g���8�;���@�W=Vw��-���0�4̦Y�/A�˕�"����zm��vٔ���f���'��nx���~ȡs�>�Eב6~��YZU�)�4�2�_.8�@���;B��5u��ڂ�"��WS�tmT�K��)���9{/˔�c{y�-Ƀ������h�+��	[�5��z/��9):�׈O��>:XKorr6O��3�@16 W�mU��#�*ĵ��:8Q�2|B|�Y.�Gx�M}��t�إ���/K�0q�r�v��ңU�5��tx�!����S��)8���gI�!�5��iH}f�oG-��o]2���8!6��e� (<�f�TI񔀳�<hƠ�G�q�h�&�ԑ�2ų����ϽC�d�6�K�͕��ey��iM ~̵ኯ}�^{3$�
qpᷠ�c(ț�������.�d�7܃����78מl�S��x��C�&����T�r�I�
�My.�W[s캃Z
LХ�J��ga�zW�/v.�Ea�~|�z+�ښF����C��:�B�r3��):yjx�a��e��ܘR9��Y�`���&S s��,��HqA��*{K>��3�P��y��1�	��:���`z���]���יӎ,J�O��@�����M&:}�fۼ����e�o#l���w߱�6���:,w_���au���"'�C@{5���/���d�F�>F�/�gy�ؙ�w�����"����q䮲����w�H�j��.�Dm��~�Y����ɛ�NӸ��F?Ē�����N����A�ք�LJ�w�/�ʁhz7�����y������v8�_���򕰽��7��s))���ߵ��)t�&���̞ƪ_�rǫs�~N���׈J9��ŏ�E�"�9b�}���p�����a:?�*�р?A�M��]~�wS��L��&m�-�No��8���pm��{�=-�*�`����iKw6,y��a������/����e�?��֟r�CZ v��oc���YS(�M�`)~	iT��@���Y�4���9#�j�N�7���%G� ��r����]��l;ZD�B\.�:��/�\�Xs1E,/g�"hZ�������7`���=^ѓ�6��ܞ�,��y��SoA��y���ˮt/�{n��@-����1���ݬ:c��V�^�P!>��a��ET�db�s \Xz�{�ƺP����L�8vg��^����R��z8LK�h�����|�V��|'�H���怏�╌��g��N�m8N&>�^B�\ Vu�=	I�����|��c�/;M
eDd�kM"��*_����� �g��m�x�υL���D��nF�xQ�m���PW�m� 5��A�x�K�3����x�� �Ue��sUE1a.�],��Mp���8i���$G�}(��F~�i��ut}�p���2W��c����Hٮc��E�_g6���t���p�gؐf�r���q�y�{�1������Z=w�9ͬ�fc{"8��T�|{i���uer�C�uO@5e@�mǶ�d��`����4!T H�N�9����x��N�	-lM��"��X~�ie��5���� ��x;������X�8� ��;�s�Ù�n��L�r���K���)g����{ �c�|�
a)~�R�٠;8��|��V��Ge�G�X[pS�KA'
��^�1й������(\eW��k�P�.�׈��ܘ�^縴#im���U?ޙDP2D��S����g6�_�;#��G���-�L�M1��"�u���HQ���]i#�ro�J�/{p\v�g3&GA��Qّ�`Ar��Djۍ��e+���;�4�Q~ũd��3��%�f6���a%��K��U��)��2΀�GQ`�p԰���<K�Ns*/�\Cu��OYѠ��:�@^��%�OE��&:"p�F��>�o�/D�iG{�T�z�k�Q��F�l��}�)�j%]�7��ס%�5��`ײ��ty�*ҥ�[F1���껤��2n#�H�w�c��#���rx� ��o��%�Ή0]��9ĳαu�>.ˋd �B���Ny����gwE��:/)+���Y�ƥ���ߦM*�e,nў1y_k�j��2�������d�jS��[7��]u�;23OrCm�_��R���Q�DEeu����"�{�گ�.jRj������'�[p���A�(E\Уj
�����\-.W*��נeI�t�����BF�����59�)�~�x
���R�ŝ�6��~���2�(�*���Ejp'�U��x�~<���lP3�#,����C�ݪ�c�f�D��$,�P����U{�.�����߶.s�|�`���e7�h�v07>���l���Q��`�B��j��Ai��,����ˤR�>0XAԗ{ ��a���_ޓ;t�a�y�·�P2Mt�&N��l�<��C��mʩ�R��q$Wc:m@�FAc��v�OOQ�@�lb�%�1ѵ�r������jߝ�lJ��B��u���1��A1#S�`����Ӷ�pYe07o��3۱5p��iZ��W�0������㭝Y�m�1��/��������q�"K���8�z��$ˋհL��}�>E�ҏ�g'�ŁP'��Nb����T��~>$*����-�x`��!`՗?:d�޺0�ѳ�ȤNU�.O)�:��_�_�{��4Ӛ����w�Oqތ��Z��=�x��M���;H7!���bxc6�����yƣ�e��
��&�稷��7�|�	��76ݨA�>�ݽtj�uA�H��3Fq��;�����F&NQ߬#�`q����);e�`�G\[4�P�l�g$�gQ��oӚ����6�nZ\�o�5����_R�b5$!B9��x�ge���,iH��0ɱ�i��#���L�Ӊa��$}��g�+����ƄK��� ��0S&���{3��j�x��-��I}��әʁ���G�
�����i}����n���M�?�;��XM��M���R��ǀ�4R,��K $�������N�[p ����NK�ts|���$0R��3�?j�c�^˿gS��T��>�!��ۙ�(/c��].,NY�g���������u�`B����*����K����}�i�Ue���h\���E0�W"�`�c�?R��Ա���<����l�[�q�B	U���,���J�$��Y@ ��%��	��^^,b�A����f��z��h��<"g����WU��oM
xE�5��
��\ ��4�H��h6�`�O���`��])����G�?�ȠQ���������}���޿v��3�����X�HԔ�4��πx�qWx�]M/�V��>L89^�lMt��M��m�P �K���u{$Q�H�tԉIB���o�P�ˈ5�����-�N�M>�^�,�b��M.���*�F�.	4EA<'�#U��Vzg�

@i؂�%��M��&�y������)]<Ϝ���(��0ai�ʀؾ����/�t�c̠IFPc��W�]P<��cj²�ݍ/������Rd/+�9�{�%��l9*0��#;�
���>4PrŅ<oZ�Di�M���"췃�vha������a��7b\�:Y�'j��;�$yB+_�a)^a*ܝAc/z������`18�0x_��w2d)9����$M7S�ã6]���lf�c�L1�|�n[�G���O�U��up�5y�HێէeUkY�+H<�N��ۛ�f,"����'���2�oGlŊ�,��w҅�<����v�ZfR�_��b���/���&�b�d_,�ذ%^!�>@���A������&�#c����E�����</c�sl�э���FfA�v�K$)�V�B摼q� �>>�e�ɇk�C�/�}�6<�љx��&����u˷C��8�����k�i��6���P���%v�K�]�윝ycn��f+�έ�;�+s6q��V*�rC�w�Y�w�/@ �?2%��9����2\�A\H"�]I?�Z�^�G�*��T�Pv��1@Xb�K8��~�xR�㲆,��]�d#lX#��؈5&('�T����e��rO��̖@E��O֯K���7�9��,��k��P��R�{k�o�%��T�� �9�.�;�$>MEY�b�/`���Qsj=)��"	�$a�2f�8Q�5Kq\M<�Oi��	����P�Ul<��R'r��?1V��5���r��]���Tl5^H�����|]�Y0�vr��_Ͻ��o'|�������z��i�:~a�%�Ok��c\|�cC���S�쪔��d��r�0ڀ/�r��'Ld�r/��N�ht�L�ю+#�r �3l+%C��G��H=X���	-I��������uޫ"��Y��ZW��i�4���P�L+�8 �%~�fR�R�����4��`eW��I�_$~��]�eP�T��<H����xP�߉���GP&xo �0���õl+�Ӵ��A��AZG�C\H�{]�Y��  �7$w�i�L�?:�Y�*~��:ш��9<J:�\
�R��B�g�SKv.��K�Km����Fa���R]��G�>r0>�A�M�!�Ϭ"	��Uv��AE���r	`�A�H'7�]�L8���t(btS����PUA�$L��|�`�9�Fq���6Z֗��zE-�᛻��m�����]|��)��Ծ��Z�0���g��v'�W�m] (ۉИ��D��q@���D���"����xY+S�����u��:xhƵ�K�ؐ�b]
��1�4�E�m.(v���ɇF@��>�K�2�N1_+)�7�<˳�99+�$����W��Jt��p������?k~Lq:��w�!���S��|j���Rn��zx[��}��m�0,/�Eb�(��u�{�6��~'γ��&�����2��A���Y�$F��B�Y�F�C�şC�P��D�C�� ���aV�I5�1��9
i{.��yԮj4x��K��-amb������y$���(U��ù�Q �C5�����y9��t�� ��w�x4����W�I#���\	�o�U���;�����{���?k�4�&�=�۽$��m�ƈ��	��M�V���tU!���i����Ko����l[�����=21>���R������<
��KN&�ο�iy�Yc]{� �M5諨��7��ȸ����ı�죮4_h_��#��:��� �\���Y���T�B��>"6�����I�a$VQ�D1} �W'�סp���۟�y��fĦ	��A� �ʨ`���*�L����t<����C�����H�o������4c�]#<ſ�$w�ԯ��@�pE:��Ǟh�G�ƾ%��dZc�����#_O�(�2��W�b<<�ΠJX�����9P���j��4�sa�� ���:k�r��Wr��Z���5r�w{/'uH���� ���ѕz�������n�d��I?*COO���k,]�.�`
���OE�U����;ҐY@��>�#��/� ]ZX��B��i2�\�d�6�����UPR֖�*����N����@h��zkX���V��8�V����.�ڏ<X���	���Ԩ(��f�� ���T��,iO����#?����V��~[�J�G5;2|u���5�2��I�(��ދ��.��M��ְ�SO��ꌶ�f�i&]<ՓZ�&9�h@�l��N���ќanp��!���_<`avO�څ*�������T�+&����J�\=���S)U��vd�1kc�*��s!^q;��OU}��"�B��)-��(bt'^cd�r���՛C�і��n�؆�����2n�yG�P�܊+�b6�,o�0
Z'$fn)���Nu��ΰ�'�˵g�4p�(q�g�����r�ܖύ9���z��$
1��;e����sYAŷ�hF���ez`�l�Rj;��9q��$K�0ld7ΰ'4�c�J?7L���_p�g�{�^=r��l��G����l�I�,b�g��&����<�q���s��?��X�nc�>�(�'<��dt��wg�M�$A��C�Ty� 2�h#��M��CkR��[��I$� 
=wv䃯ȹ�~�����}V��9�Dغ����{K�o��s�\/t���,���vY�.ؐ��1@cSCy5!9�E��ب�:����iM.���Цv��X�#Q�~E���`I#d�6���!v���EV<����$`�#)ޚj�W����N�꥟{v�݈l���5�C:��:S�("��I�����=��DΙ�N����)_�4��/	b1{����W�E��;
<�Ӫ.�1�}���������(<N�������c�2��+���_	��0��	���M:r�*�=�27���^���3�=�(������y3W���Jn2$0%��u��o���BF��ЙDv�ܖ�(?Eux,��7��<�^����Hu���������k�]mM�C����̸Ĺ�b"�4�l�o�'�|H2#4�l�Y]����++^�c��_>�9QLB���_f	:��b:����5sU�^� ��4��`@�j��c����8���pߥF��<E1#�w��OQGd6�ڴ��c}���ui��"h��E>~L&L��-eN��p^�C��L����M�|�l�{�ys�7+�4����a�{耏&��k=��Oe�i$��U�X�y�7�����T�.��u���3v�� m�yYz��[�,�G3���s�!V~r#��JlA�9�9���nr�쵏ܙ 92)����D�|�S%��{��4R��?��TퟗZ�}���uUO_�e]��+�5ݑ�jY$P�}�&��o\(�#e+��7S�����;��M[��í �s~�˟
���k�&����N`}:��:~s���,�����5��م 3s��W��hQ��[�,�k�C�߆���.yG������	�)�8��G�1�`14G%��� �8��r��̉�:}�;t�a6��y���l~��E�f�#+!��ܷ�^`ͣ��͡=���u��+o%����5�,g`���=�C�F����x��q�)��\Sr�����]��������� �6��`Kv�Za����$f=]��y���L�œ��.
+r�=����u=��$ȎM�7G��tu�\�ѓ���O���Au�(`�p]�a1��3-�����q���Qgm�9:=oIr6x��F�DE�ī§`�K��TY�W�eYX�\� ���o�t���V�o��.���d��ɫ35���9��E�+O���P딹�X:���@�$��z��!'o}� ��S�_��9�`��2oG��&m � 0O�kk�[,+3��5mZU.ciV���������� �Q���ڊ�n���k�퍆��W3*p�h���@�U����A�z�Nz@"����џrB선����ݢ�_rڙ=��(d�R�@�ZRZ+Q���U������`�:�^Qx��쮟P�J��h@z�CK`��N��^UUY������1HX�����g+͌�":T�b���朕t�g����H1yX7��;F���҇6����j���HT�/^�\B��tM]��"��m�����1��Ht�U�Ϸ5�P��Bz&\����+דsc���n�}�qGo�e�����*B<\Ǯ�Ud�Β 1_�t@/FU�5�X(<H���C�z�$�^(��9��H 흮��F�L)34"����#�X�4k Ƈh��f_S����R霱�4�A�-X���񄄚��\�p��bv;b�l}��z�p�T��v���M�����/^��q��k�N�k�|d����N��@RETO�-�6{6�y��ț��D��\��3�&>
Ej�d�GD]�(�Ī64��_�/'ecFOġ�C7��W����/�{)0�ͷj��Pɰ���,A����J��	�ԃw�Ӯ���e�P�1lT@s�b��p���?B��������6o,
r��P����G-u��F��*\��eF4i3}oο>�iy.>�;���t���7�t�����&���ʰ��Z+���U�]H�nSyĉ�55AuR�WLx���C��m\:��]��e�A���;�[�3�� �_�of���w�m�!>9�KB�Ѝ��Yyk���C����5��V��k*E�k4���Kp�1So��V#����B;W^M���Q�NV�ի���3�t����h����~tʸ��:]'K�C.�_K(&������	�5]E��ތ��k�v��&$j%�Ojq6�t�����q��Qo�>����bL��i�m{
��Cn3��eC��~�h�������f�UG)&���3R=�b4	�ʖA�cl�
@�C�59I�7|"J��
W����lzgm£�����=�4K"9b�����6��f%5�=���(�j��)1c!�YU���4�1"��}���Z��$[���>����o\�3����Y��� ���5�O��]��.#���I �4���0,�;���j�����zɣݯ��Tg�t�t��^F�@X<�[,$�?R�F|J��B�~��#�>׳G�ƭ�gF ��q���|�x��5��k~��G����!yW�t�^Ә��ۦҭ��~�#8j���8Zɑ�a�)�o����H��'�!x.M$�?ՠ��hǰ�GR��S����?#$�Edґ��-Xg�`�&��d��ck�wCb�/Ƴo$��b)�#�}1�P�j�����j����b����lܧ�2o��p�3_��Ruu��S�A�����{ 3-�_��lP�6�L�V�>��iQ0�o��Y0�*$ذ�f#4y�4��O��|�`(�!b�MOʵa������+�w����X j�J���&�Gr_�Mȼ5�)����yv=2Ceݳ�S���&��Z�oltݜ�>�]����J����/���֯8t��vD�6mq����d�X� �+��C�1�Rg{�:���O ���B�$�Jx�%7߀��Og5�c�̈́��6��#x�;V!���?/�������
�z}�Ŵ�6�Ē�_��*���B�gڠ�/WA���u��T�A@�H �%�+���p��{Ԫ��-��9�J�)_F�"���m��v���m
1�6"�3d���+�S�W�E[H�7�\b#uп�L
$��i,y=N�&|���+�(�7`���%��]!د~����>������W�]hym��؞� `������MM�}�����ף�@��>�k]�8Gn:l��e���Vhv�.���L����
_�튂':��`�wD����OvĀ�wn��.xj���W+���Y����N��W��?��l��t��y0���<��.�f;ap뛨Q���9K}��ì���aL��w�m,��р���̺pD�K5�h�=d������ ��@#����di/���$�^��g�eh9�ں������t�ٟ�#=���1�V�9)�������Um�OHSj�r�����pE��/���	;R_��,�H:y��Y8!����!uA���|�c)�2��؀��b�I�MB��A��T}4���^�M_�#��ÃIA����' P�D�&+O���E]��%�{S�"�x*�LɆ�oR)vL�D�7Nz��^��/'��U���yn�r�hop=�тM� ��>xX;��b]Tͨ�Yr	�?B拻Z�����e3����`�w���7/�>��Lyа�s����aTm��]�&�r4r	.����\'E8���8��<�vS�G��F̱m�k������H����K���A�T���{ޠ��G�����CϿ��"��]#�V�G9���*5�Pybz�)�p) ���9����:E��؄�V���!6�r(i�����~�{V�!�2�s�%���S���{�ԝ���H�9p�8��Wb��'	�dԢ��������>F�)I �b:v��ڃj-Q��M8�lH�aJ@�j@���������q�����-�K<��Y�̕�{UqZ�����[��Ys� w���J��b|��I�0Ħ0�Y��� e@xA͝�ZѲ�$��G�φ17�1Z�On�6��!��K�o�N�(炋��[�3\� &eB���i���5�V�`K�b�s$ߏ1	u;S\N���/�-	d�&��K!|3��������d�����t�����rQ��-oX�ɚ��`�	�7��n	/��*Gʣ�05�K�76T|i�%�T�u:N��M�Iu�h�-�+�� ���+��^R�n���R������Q������:�y�tz�!�,�oX���t&1"��7R@�i����f ��3�0���&�q��n��QS.ʝ�m�v)��#�����z���~��EX]*���~��LV��P`i~h}��l��5F�M���>��z�s�����c:9���eŉ�諦J���s�8�ht	�d����bL���&黰��w�;��*�b���^��˘���t].�RA��Fx4-ea3�nWQ�����d��� 7�Dq�@��Q5�.����+��'��<�_}@#��곕 E)�,ugG�b�f���$��๴�96І=�.�|]t�:-3��(��V���.�5T��n
6�9���꾤����i���@|f}�J����5���:���o\��fG�����I�.�c���H�*cݤaz49�]K;F���}�d�GRU*�u�Ns#�c=��e�ֱ�RO RIF�_�9��)����&c�Z�C���J�V>��8��5�z9��o/���>�z�E~v����M�|	V)��8=��X�`�/�>r�v<֢���d����b�l�5KQ%񁙺L��Sn��'8'T�,�	"��=3P�|,�p��D&~�����M�
l�y~�oA�I����F%�2�x�>O���ػ�q����83�dA����t��f�Q�Om�D�m���$�L�c�f��:Ykꟍ��IЀ*
����C���N;>��G{�L>\/1C�V�x-��B�YI�*�������g��h�X��5�-O�9�:t�"�@ў���y������X?�e�|���g;�����6,%��I�z�L�l��ۺ��2D�Qߍ(vҖ�1_d���%q�IW�0����Av��Z`�}Lv�	ň�G�l�ދ׭�
U�Y;�X"^���c�B�:}+�5�\$���̛K�@4�pAC��i���P��Z��R��2V
�X��ST(�s� y�#�����9�VO�K>L
�F!�"�G��CPf^06k�*�k%�/WZ
�P�?�@8gCEЅ3�$�OD�;vzߝ?C�hF��aXr�.�Oŉi�Q��E�r��,%L���lr�]���s��k/� �����&Z��O<�Tx�[Zy�w� ��~���������NV�����]���Fb��5�Pܸ�YJ���������m����a䮮���������g
���l ��Z���"Z[&ت�+t�Qr�ƌ��4�D�d��x���Q�Uh�z{x���th(6$��A�����ɖȫ��[7�hC���q����wRC��P�D?����+��C~�irGyĂ@�⓸B�&��NT?lxǎ��> �<O��	�16�1�|�Fl��=����-�ȧ�c���%˰@�)��?��A8���WʸW�N�!�����Nc�I�?w���{ЦGӖ������ۼ��YEս>�@V �w۷S4�}(�qa}1�Wt%b8�����x�,�'\\�4��+J`$AZ!V��ك�C-�{A0u��;/U^;��p�4G<*���<7化�(.�t���I=���(��z�M���u�-����h~j�=L���Y#:?��pUa�� �����nsa���u����[/�N�M���+�`QG��w����KF��N,�z�����Ǵ��׌�\=�%]���Ie�2W�q���f��S+��ǝM�`���]��QH���7��ER�JI<*�P�2y)E3�^ǉ�U<�|h#G�_�aD�S��?BU�[4I�*{�쨾��v��Sgoї��4�@�:JCЋ�/3S؜7��9M�{���l۞�֞m�0�߸!7�>-fX�EA���R=��a�Zע��G�7\�+L��Xy1v�]c�:4GH�8P/�ą���E���(��|�yQ�w�:K�r��1��s�vV^P({YZ�X�䵩Dol�k)% ����R9�L7ky�ò��W�+��Q8��e3�Q=Hv�}K&�JI�25c���L$�i�`�ͥ���^�o&�*Lf�	"�,N��dF��q�t����[�8٣$��+��r.���ԑ=!�xþ��3���SMF8^�D�� �%Q;��I^S*�������o\/R���P^�ϩ��/�X���K#xLVA��+ԧ�ի:����M1�GO�Y������h�{�B��/�C��-���������G��n�d��v��i)Pv≦H}XZ$ҫK8&v�]ف2��Q�S9��C+Q��G)�O~�r_6�ߛ
1��OC�`^����{_��F=�u�G�$r'F�9�����4���_�@�~�m9�".�W�A`mit�8X��8���^X�/�Yc�0\���U���X�/�U�QR���{s 4Ո��#��c�vH���U�Ao/ΙU�h|��j3ΥX�`y�9UH�q�q��G�щ��R�)`�"{��M���f�s齃��fg8o�x�H٤8<����7���[}NEŉ�I �l2�Lܢ�(����Z1��2UqnqIj��ۏ��d�r�шg�zP���э���t���B�P`u���Śb/��U�G
���	?H/�쾘~t*Q ~��F�6@l�yb�*�>w DM2�˵�We�قU$�Gyh)ehmW�i��"��|[��N݁�P�rQzh���gެڸ]-Bz���וo��B�TX	�p���x���m�*��2Z��S�ؗ�h`�o�KeH5֛�^�ܦ�u�o�H!���]��t���(ܾ@��Q��W$�������.��Ty���Q�X�_�ou��H��a݃�
Z�6����Tv5�/^��=��Y�$�R�{[����w��FYy74֎L��=�b��-�\�?WK�%!IZ��m�RIh}c�_�FW<?�Y�׻����s5���ʝ|�wԻ��O�EEJ=��w�Q,��'��u�i�q�����+&�1(��|YlWr���w�hY��k�����v�cҩ�aa4�O�Ry�ڋ��t(�P4���ꇁj`CV�f햡cV��|0`�}�"���z kP�NpL*'{��)٪�T��=&`]
��d����*P�m�C�r��j``�Y�n\ח�00S�c�Ye,lL��n��ۉSp�� =X�?r�&�{\����;�0QfR�61Cc�Dxm�
���bt-i�ϫ4y����b�ԋS��(L�
���\�}�9�M��� knf�h!�Һ:�R�. �I�%볕�?=�Y�l����e2a��!?ys��;W��Hz�X�*�L`�)�OB�oR(�W$E ����4��Le{�-/�^��l�6j�L��^��ǹ�@..���X�6#�)8�#��q���xX�a��hļ�N�f���Vu���%_f�oM1��Z� |�E0�m�T��̇ؗ�P�X;W�6��Q�1��Ճ����w�gV
��,`��{C�T�$�+U�G��Z�P��x$>P��\�������8�8W2S���PRIg/�6;�7��
�Yd��?���C�
K���b��ӱM!�{��<t�9��9�]N������J�S�X��I�#���R�5n��$��h^�1�1Gk�t ǔ����Z�Eh�� ��n��%KJ�K��;�2��o��u�PtnMW">)�x�H`_�Q�ɞNd��.�`n�^�:�]���it�T��وn�hẒ�	�R�ݩ�~ 9C�n{�PI��ςV�+��8sه2� ݢ2�:�`+:�L�0��?p˒�#���P���ވ
6_թֺNCG�v��s%�W����8��ˑ�������_�۸���/��y�j��c��1	zao.�i5��NQ
��k�D������,���M�,V�ȗWN�7?�&��;nIP�Y/�/_�����w��m~FT�$�0D ԭ�F�,Z�w���ivy8D��������^�ІV��
&��C9����`�eI�jmQ�N�,;6�*K�	�x��M�t;�ۏ��l�I3I�#��l�04<�*�p�ޏq�e_e��;4{�/�Ѧ=���g�:=Y�j\��Zʛ�	� /*O��7��R�	���:�c���z^
�;���ko6���6a�{��/V��>����b����X��ʆ�e���a���I�c.��S��ae½fg`��˫��X�L��:a�,c�ai�0��>Z��K������t�B��F��9�$HЄ�̔*��ĕь�h�:m2$+b,3U�m�@'�W����
�r,`�����D��Qc"��vJ����DE1�Ɩ��[՟`�����=>F��]2c���0�y�31͛nH��(�JՕ���0싅�BP8M��y}(P�~��ʒ�ˇ���]]u26M�Xsă��>�hAВO۵4]�U!��c����X@��#%�ǩ�N(�3I���2$R4~5q9��򤃍|t'�l ש�e\��_���U&�׆�U��י�6�hQ2<_v�f�,�u��^��ȴ3E�W��Q�Pu�8nT��U����]G��G�V�§���ʡq�5;��
�[���]6e^�ΌN^���!7���������vb�ȷT����n�ڂ��L����n7�5�K�]_5�����1�~�@�����(e�D���O¼D�9P�q�Dm�@J�ر��b�YpNޑ%W��|�1��eN�d��?NM�{�>�vV#T��b(��=ƨ���&r����$~8�P��9��Ç�8�Y�P����g����v��P���%g�~p�ѬT-�[��޷:�\Q�e���?F7��C7gq$�q�t7�kcit�BFu3ƒ�4iw�,��M��$V�Fl�[���d5G��Q��{pH�ޣ,�щ����P}AM=Yc%�d�ۥ�~��Ka���a��d	n�GX$̚�/Ll=�+��E0$n��A�|���n�-k�ߩ�����>���׷��C[Ցw���n��:Rd�4s��ry�+�x������5d$ť��w�	�R%�:Ǽ�q2�xk���Ӽm��/@��b����1E���ȁ]X�&�����`/dfԭ:U�v������<�TI�fH$��Q�ϳ��b�$͠
��I����zX�o�iO��z���ᝧ�:�PO���Wܡ#���Ӟ��h�C%�L����<�@�b4��h�}~8�NJ�C\���!����Q��t��T�����Ɇ#MP|�ѵI���
�X��Vņn	�aW6Q] 7�c:S�(����M�?�כ�Y�1F5S��]~50��eGO��S�H�X����A_H�5���.<�f��H+Q���b�y� ������5�&��Pe�����ZR���)A>��bHg'%�E�	�ǁd3��B�iN~L��sx� �&ڴ���JL�b���ЇM� %���8��x����K�V���xPT��\?�~Ru��k�#���j#�ݖׁ9H�Ku>��k�(����{+@b'X%�xD����'(���`�1�u���!82G��U9gkr�I�5��5�[�� 5�
k�VU�wS�@������ґ�N�b���[��w�l���:7���V�w��;��#�~:~5��{�_��}���������fx�9�M=����{o����BG��t��D��Lq.hN���%i|����M�C�PLY"�9�+��9n�֮8I9F������"šv_|������_���M�hK`��%ZQ�W�Q�;�%�U�hGGR��Y���W}ŉ6(��N� ���:WW�j�s ��'9;�o�m3A�)%*9d���� V9��5pJ'���~Z���J������@M��:���"0�[:��J�E��׏��S��b�;f���H՜�� v���u�� p\�$3�isP�,ՓYj��>�0ǧ���2��J*<��ZB�
+m�����U�	�L�+ٜ!��z(_�Er\�~�W7_��b�a�b�;O�Ƭߍ�	j��hlq{+��j7�w)�h�k��^��CJ��D�q�B�.w��V��#�6!7��/����S��)����r��H�M�[�F�"į�o�_���Of�1ٰ����0z�o�~�D���A�i�g��I/j��rF�n�K ��:�#\�R����Bel�f#�>H�PK)��"g7lclz�
�1�~9e��~2�ߟ�uT�8�G��E��Hf�YS۪w�
���.��U��4)B��9��h���6��P���
�ezf�g�$c�Ȧ�����R@�.�9U�#��@G& W ��ߗ9�Di�A��yd[�A*hԆ�����	�#Ҹ��@'m]�KR�����	r����=�&�3,T��J1/qg����)���5��� ��0���ט���߹�	''�n�-tbא�(�.�ǲ�-_ڣ�g�����'�1)=�WI�p\\�ǭh!��;jv����ս*�FT��+��CP���ヴؑ9��N)��&0c(+��ai*��tr���)�Dƣ��F��xd��[�"o�V,�d ��˛eI9�$	D�*���P	���ǔ�y��
k5��٤���O�SO6�~�!Ի~���P"�oc�\��iS��*�f�5�x��U7bpH���C;
w���X�m�?!ͤ���ӵ�rD�<m�����6���y ���B��뜥&���rj���C�Qzǵ)5�Um�B���O������9v��ڮ�{��8Һ�|������8�8ҿ.�=N�CfD�ށ�y ��;���+���?�P�X�����ɒWN�^���*|�X�K�mq�I%�p,�yt�5DF��/\��.�OV̥!���	�����%H�����Z�R*\�g_8�i�,*�Mk�	�BA��k��"�	��ٜ�.@+}�+�mk32�򚥗Ф�*�Xa�o��Uߜ��CH@�KM%�P���X������<#����&�U��5���w;�ŷ�h ��}�韭���pN>�J�e\�P���^���.��%���1������5*B�!�"M[؋W�C�aq���
`��(MT�������Ů��F�X~0b�dq�-���ۄ�~��:�qۋ��+^��'�k�'d|�=.�E��L&�q�$���t�Qf]ڥ6^��(��Ёa��Ê(�޺����+Idt�E��[F�v:�[�Y̤Z��#X�,�/�v�����=�--�Ʉʷ��UM&bZ�R(���ŔO���IG�X�n~4Kr�ğ��,��J,mL{���мIsWD��4�e���ܖ���f�eH���T�N��{���`��}�CP`��e5��dtI0@�;�kγ~�(5@CZ@m�XM��<f��0A��<K�u���������\��z�9�8�2���	�������I4w�캛O׺(V;��x*E�)�!��9��رg�!+ّ�"LJ�I=����3���[����X'�
ng�ӛ��2�/BI�{j�9�p��5W��^ݟDYʂJ��P��@C�+�08��į���fS9e�L�� ��7��z2�.c�n�Ǡ�L{� ��`���(Ǽ��ܖ�n�B�w��9��"dbylܶ9��Q���I��Cb.v��8�<�4آ?9w�p�$ Ͻ}6'�Gv����A|��0rC8�)�=������2�]���9+E����z��M�M�-r�M�T�^�y�ȩ���~y���ύ �L�.�6.t�1yh/b��IMr�%� �$�1=�?ą�~b�n�炋8�1P(DX�#a�^�����4@�t�hZ|:�nCm!%�Z�\z�ךo0�
�y�P(.%��p16�ƺ.���0�gul��z���%��Ǝ�[������5|�_4IX��3�LNoZT�P���a ��5��槜�����]��n�u�<(��vN�����EI8d��Ywd�����˯J�$��0�g&2�!ڟ��O�k#��~pD���YI�eV���
$���=�b��Q���+�
Vc����A�H�1b�����<�4��1ލp��'���lH��"|Խ�`:�_�5�=w�x��!��xh5�R*�E�޲͘Y��,[�D�=�h��p�_����3������p�1�&��-.T��=��.�o�>w�>���y�������Q"���x4ǰ#���o�����&�#"N�<����D*)�Օl�7��g�椌Ω�{r���6���xm����K����O"A<x�C�X��j��7��-iL1���R��Ku{0py0�u:���@%��)+�[���+z�w�NG�{d�Iп����(����ʟm���~��w� �𲵻�ތ�U ��A2������2���ia'�XO��n�C{�I��-��!�ƃ�b�7k�.9�l�b44��K@3��F����PB���rQ�vO�?>7���)�M(�ax�|�+2�/=���X-�TXܪ��Nڃ~����ى���PY���t���|�5���*P�5X9��T�VF����/!��xE�(�(N��F,(�Í0��]���
m�d*0�y"A��� k&K��;�CIp��#��+�u�K�=N�i�M5)��Ջ���\eJ1�3�<�_�
���8[�-��>����h#����;�#L��I?2g�!#��M)�:9�%��q9�S#H��U�\��A�bo�ك��{��zb��������bN�y���U�q���/A�G���5��.0�9,�~4n�h�mM�0�nt�x�-1J��-�%c~ڎ�l5ΆJ:�a�M��u��m�f�PC�o���S��.gQ�	�S���1���KؽC!bO���/��4S�3��z�C�h�vN@�{ Zֳ�.�2=q@���Γ�{��Yݭg��I��?�D�[�R��q�j�ڵ�ڏ��`g��m����u����Uxl�����pW5�;����Xm�A�n�r��գ��*,�8�6�$qk3{,�y,���ē��Z���*�K�Ydo�Q�I�!٤�[��3��\9?0�N�B�~���T˫�5xM����ct�Q�׶x�E.D��H��,���c��nz�� �ѭ�N�(�����[o�NVLq�'5������{����]1f�.D���#D#K��|���GG��p��T�$�O�^�Q�i�f��0[��hC�F��g�SZe��K���y����.�f�G�67�`o>�
ڽ�{��t&�4�k�mיP�T��G!������*ה����,9�wuF�����GZ𗶸�Y�E�dq'�>�L�V�UA�w!j��'���P0\Y�uj �fR��,�nB8h�����8@=ؾUݴ`	��^ݧ</�}��*��|�/�ĶՕ���X珒*@�11HV˓�,8�g�"�,�9���KQJԤ1��񎄷t�c���-� ;g��!�����I=ve�ᅚ�wڳ�ղi©���Im8�`'���2k�H�d�(l�TǘVB�l�2��C�F�E�?=�	N�W�U��"7P�Sw���`tΘ04���Bv���j��Gq;��{��s:zx�j V�B,2�8�Mޱ���*m�\�#nF-�r������қ/�;�Z���_&EP�� ��xH�2a0>�;nr����0j�
���1:;���d+���~�ǲ�]U-����M�!��p�6`,'ג&��5�R�nf��I�sN� �c�o��oJL�-���M���7��PIV�>Z�d2��Hy@�MsC ���2@X�k�A)B@ҍ/��?RD�%_��¦Y��"�k?��Y5�a��a�,������K�]�kB�tB=��y��~�1*�Ԉ���� �;���L#Q)�E0���8�3r�:'���zU�&��%�U��*6��Y�?�)�5�W�n�C/;x�U���&�]���C�[�Oz�39dO���ãy�:�YW:����������PEC&�]�y4q�ʷJ��#�v�jk����g! ��>]��v9��&B�d�/f�
ӿ�5�("ߧK����\�c����- M�?i�s�.��/!�A�˱�'E�-��H�E�z��������wLB�dl쥒^F�q͎wm��/Z���<���M�Tʁ�Y��y��v0]�U�,��R�E��΍{���7`Ԟ+¨[Y1|�׳��YH�T�/v/�\����x�u>�n>�C+�+?�QV2!�VYS�v�, zh8�f���������&���jH��%j7��:b14D,pM�\����%����Ҋ��X���wVG���U.���	�v1�y`)Q�g����h�ԌS0i���GL�����j�\8�ie�P	6�!K��q{p��:�xY���&Qg+�ձ$�r	L��
�A����r��&�O.ɝ�$�(�ORO�z&�Pl�A�P6��
^|�	���q`�4������e��|�0�uf3��g�EnS��^y6�ї5��\*�Ã��`�����g�����n�_uY��F�
�9�N �}ݱ�U�E������^?��n>��5��T���Σɽ�I&��1<Fn�I`�_^�ؘu�|���RqنIw#+?���P����N�3Ed��^]d�>�A�&$��P�)��O��q�3������!�$ ��u�p-���&�elJ]!?�����2	� ���!a�7��}��.l�we���<�w�R�$�T��+)�: ��n����b�'u��3A�)TI��}�Ǌ�tX��&�o=S:���	M:�%�Ѡ3���>�^*3�ɯ~������6A#0��������R���)Q.�q��XJ���m�a4KW�Q�a����f}f��CLj�T�{7A��f��<��� �$�I(2�Q��p�����U]U��I��$�e*~rF�Z@Af����h���N��p�������m�O�,4�!�Jµ��j��������4|�jQ
g�1��5-��}x{�5���1�\��:�"��j:��`��iw�%EΣ]UZ���פ��N�t�G��P6H�Y�sEA8��,�����	>a�uHćt�luƉ�e/�i�0��� x#.�'���I��~[x�w���v6|�|��r���<�μr�{�c@YX���uv�5��s_z&�L2���_]ց�8'
#Ts�lv��Yh$�Κe��V[�|����9}���^$%�]-/�)�+��/\�&��s��]Osq�x ��U�]^� c�,��ENqY+�P�`)a���N�I"�5'/�f��l��}pV�P�)P9vgc�!����Tc��v	єqj.��g��I���<���@���R�"�k�����Q��	Q뢲/���^��<5�>�<>/�����ԣVW�,�>3�*fl{��G(��kuØj�}�U:%X�7J���N�����؁�*�eQg�?˰��F�
��a
�4�;c*B*� 1�݇��qI�o������5�eq�d�C�_P\������֩���G�Q`��so�����9�Rs�ZdN8�G�}�[=O�U�p �d�8�?�es�/yi4~�R7��Z�Cr�I��$j^J2wb��7�}�,W�px�����&T�s���"̹�o��X������֙ǆ: #���Q~�ٞs���,��7.0�$�F+oW�,esf1����eJ�+$��$�۩�<�|Ȑ#�t���j�ok�ýf!�Oi�r�-z4��2�ؼ�dV'26o���S[&�,�vv�|j���JN"i�hܑsr��MU-�[��^2C�t��}�cXZ��>�S�=Yo�:�0��$>���yZ�T,�*sh�\
_D�%˶sO�J�5�o���x9zV�J������p�k�.Q���Zd&oy�ڔ�Nu�ɓ�]~��90R���2�n�	5<�����<R�a��g�a��`�uZv{��W�
VW�Oŷ^G����x,l�J�ZKK~�L��c��P������+�ü9�sgf���:� �����_=�}����Rf���AԆd��Ͻ�����)+�f�-:����^���ǉwI=�0S}�%CJX.q��ctls�.|~�&�L�86�"�C�����5g��c0�~�%X�m�^�RC}�k�eĭ�)��fu�ދ{�x��Pf���E�T�$��wE��s�m]��n,љ�*��XM����7f�|ӂ�*��z���oO�,q�Jm�C���6Sy�����ܨ%�>�K��'�������=]�aW|X��O.a0n9�h2dU�M޼�>�:B�泯�_� ��8�F��)�{ǌˍ�\�x9Z*� �ԺY�_�57:��o@D�᳼P@��M� ��OͰ��Ͱ�&P���$�An����,
�����UM���SC�D���E���
���e%�ep����F�����'$��`f�Y���J�&��#E6��m����g�ts�)�s4�9T�M<@���NvE�1Z����"���$��"��R,���.����3-p�眠����4&vS��˦`)�N�\���)�$�O'?1�Ǎ��V� -���KIDSIQuŸ�l�^49C�<|>RmR��o�{�K��63��r�I�]M��1 ������c���O"(�3�5���y��%�͉��
�<��J�W>��m�sk^��0�'� �f��B��xȋ�V0��2��Q����iL�~G�{
�ƅ�]�2�k�DԛD^�>�r�-$P����n{��zA��9�Q	��5�,Cat�J� ���/���i[�x ��棚�'�5�$�}>
;���:2�jkY������|�wQ*l���������P�Z�����-8F�0�M!��$M.��(�(�T!�w�|2e T�:/`�1iQ]Sf�y�?N~�h�rX�~���P�%����*��|�2�֝�
�45 F����6�:����h�&�	j�TakN�r,�z�k�m�t���*���LߠK����T���mZr�QoA���c��%���CZkO.��) X�6m�������W�U�EM�Q��q�
���-WN�$#�DV���ر?5�1�r-;�q;�u�H�����=�@_N��ZZY&s�Lp�Y�J�V�b��e6�$�k�^�n=c��C>�x^�G�z�9TB��y¼Td�g^d�^F�AM<����n/Dc��sՠr����b����`+>"Ma8�°)��I%��7�kL�F��Elb��<��Ta@JJ>����(&��r_��'�$�Ag{��������}
	���X��;af�T���`�Lo����G�iL!���v�;Q�{�7�i=;������s9� H*��6Xc�W�YY�t3�ud �7R�]Q�8��A��N������U0���Y�ʮ�W��m-JudS̮�:���G�<gJo3��FGjM#Rg��wXHSǑ����)��X�]`8o�ȭ��Z,+�<du���캮M��[,�2��x���U봛rP�3���(�֙���ڬrc@θ��r�NW\����4�K��v
�qLQQK���Cu��"�<�����Q�j�c��I��!�Gӓ=0��h@#��}_w�$��V*[ȉw/��=����k���!Ga��	A7����g-(��{jH��Mf 7$ՙ��vS�h-u.��֦b��n�a��A��&�1^��?���R�Y�����y�p�{&,J���H����Q0�[��N9�����]�_(�Jm�;g�ቢ�*"���M�s�3ПS_;�.�w&~�m���I����q"v^G��6ű��,?�%���a,��*�ܑ�@r�+�'��k�
w�����l��f�@���Ԙ�evҺ�#�e����ZfձMC��B3�^}��|���"�p�Zkf���s&�зR*��Lؗ��
-���z�ѫ�{��G2��䡷�*�NS$jC��{!��/�	n�O�e6�����*���
�~�7(ֵ<���U���x�Vey��.���?9un��9��)��!XR?ċ�+�7��s�MƊ3��V|���O���:>TT����o�20�{P��mҪS�?�,#y���".�p�-|�������U�>��Y��q�i�q8���VO�v31�4����# �A��@������χ��e�v�T,���
&&�.LG�XD��kAg��������;@b8�Djg(П���A�:���%�!�?���0���~��U*��  :�P��bU~�t7h�|]���&E��*�%_�\�2v��)��ذ�bj�N��>N
�Qj�X
��ۧ����R�G�K�O�'н��Tk�dp��d#���?vn����}�)����`\ӑ(6�]uh�p�aA:'fL�1�L�����T��F�mr� ��n9R�^T����|)AW<��Jc� �B�u���n�HK������o@������e!)"yLU����X���:i�
��l.�l'~Dj��}XsRS�zE9>
z�Eצ��H��m��Jq��0L3��R�i�������+��H�IՔ^��w�qŀ�<��C��r�L�ؖ~���frlF��c ��eu����6H4�7��A։�`!''��&v9K����������'���m��w��8�� ����y�D��-���s 	���$�4�M*�7BQc9Ƭ��=� պ��;'���!�,?�u@<-Nue�&�S�I=7	���[�@?6��Y�n雔� ��b����t��~�PD/�؂#��B�v�� ��o��s��J`n���c�7!N���Ĩi��7j����*��x�|Е W�_\Α��щ�(�(��3�*e��!�A��{xߧ8� U�g���t��Q� ��TzMQ�hN4y�x�'ۭ����O�D�b/w�����(����R�a��$g9d4ﭟ[�W�
�ԅ� SDuP���#�W"j���,����*�����+2������НK6S3{�pn�u�}Dҟ�y_�]T��w��?���@
�J||���5+c��+��^��X^��G�Ѡ?�S�H�O�3�~��rI����%/�Ă�Q�]�{��є�1�I��q0v#[�ʸ��dHJo�
��� q�<|j�Щ��:��E���f�{8G|�R�((�[B�[��W�z3�s޲NP�8��� ��d ��"J���_���fo�D:����L�Y�yy�|m���K3��	���L�q\wB��+�ӿ⠟�!z�G�=������ }��闘=3�k�M)mtW�� ��n� ��l��`���
���Cn[�9�j��-�T����(�t5n����0�I���I?p|b��`��N����������1����u5�%3�e�彤C2g~.1�m�����莥�F�-��Y>��j|KZ���s���iÌ��܃芘/�{v�]�Tq�n���L��}���ϤT7�}���g)T�w��N7A��	S���2XY5�,2�/^^"{�s�q������lU����,�lįEqX��_��$��v=�q�䬗F�R��1�B1���y*2پ�ڵ�$���U������0�/>�x�:���#�u�c(l��CA�ytv�-�F��6w!���ZP�=e=L�\�?�����ע�&�Vc���Q��$ܷى��B�w�0��t@K�������"�F�
Ǉ]��4��{G�pp"���pVf����*�{�����
�P�u}�4�0��i�o!�p�Ek����Q8�p�c��5�{��duor��E�%vv��IE�g[D����F�?
+���q]����;� �����O+�je�?�e�s�j��m��h,�U�}\㍼Hu�GC��W)(9Fx�]`fF�<Մ����79�؊�}
 WO���Tx�zص��_�
�9����,��s�-P��z����KP��@!p/�����S�=5�ݾ��s���]DΛ�m��\?����_�T�%|�E�AY�l,s �X5'���q0�M�3��WZ�4F� +�$r�m�A4�=H�HI�B�s�,�(5DƮ��4������BׅE�>3=ֽׂ������h��J��e����WTc��w|$����R��7��G�v=3����w�L^e��H��=�{�}?��<"|;~�{�/�X�lt�o⓯=t*��|A;N�!�u[�I�X9��>����s+ ��f� J,���m;B��mڣ*2+O�����\,���+�T�H�k"w�nI�-��#�:�}�����)��W��:tm�˭�0�*��]3w�7����ę�c��s�2�H|o��^�R�rk�{<��
�\	\/��N�YE-Q�_0{7�=�z��� 	(%�>�6{DzLZR��;pI%�7]�qR5I�$��S��~J&*d�9&-Mz��z��;��G��g�����{w-Ϝ2�";��2Z%EZW�Z���g��M&W��0��%0�=EA�8��kv����.�t�+H��Q)�@)�K
0e��IP["r����,���m#}� {Z���жPX)֏��h�?���=m�:d]>E�My�(���i�N+�Q����$�'a�Y[��}\�O��K��~Z�	K�S�5�.~Y�nQ�<4F���7����6_ހ���~�t����)��]R�t� ���E�ͻ��ԙ�e�l�uy����e�����bO'`_ �����}�"&<O������ҫY�=�R����?I4��qM@�a_����,�D'�V�������O�}�Lb��!���~��=�ݛ#������KI*W�EV-��i⎥ �E����]�s:X�Ʃ諕DCm�E׭����"��2���>9x᭘I�g7���@J�6�ՠ;i
M?�6���H�5�M�vB�%�-��{�@�8ڙ�x��k B^m���?�˪�� ���˚���we~mo�js������ɨ���@��x�� U\�s�m��j�W`!�� .I�
2�/F�+��b�:S[���l�>�B_~��@e|汍G����V�>e��4���=���ΔV���l&�
Chӽ{=�=�ʔ��AVjF�0��f�A�P����I6'�I�	;��,����1���uu>;���n������O�qݾ_��[���-Y�����5��=�o�Gs�w�HL�����{E�u�O>�D���l�Ro�LRL�
��}F�u1��A�2z�$?�YX�%` 
�$T�ԅ�,����D�-66P ��t>HX��ި��2��mv��V�&��F>#\��Ҍ�7S�CHv$����#^�ŀC`�:_��Χ��I0/�o�Պ2 �З�}�Ȱl��;2f�x�3�,�V�#���X]ep�AUq����^�q�.�fs��X�Z/KG�I(�
��W�V��p�;�FVϋ�~q���RV�? U�l�hA�<��h�r��>׫�{���XdV_7=�����������7���f��A�Kd	��L��y�'�J5��Y�}��pG>2��x�������I�-zU}�#�hp�Ja(�|��p}�� ���V�gڀ�
�yvbB�!7Ԡ�/�v��,��0�]���M��|�%�/dWV�x9�0Jn�AI�xfZ�@�b$����;��ܽC=���~���$H�
�/~�'pw���b�����S;~-N1vz�"^A�$~G��P;�� ��ήƊ�c"i ]��o;0tc�q&�m�МI��3J�&�}�4�g��$�u�,�t���35�Lbހi�}0�{H�Dc��G=M%��֧��5�x�@k!�qq��k�j͞���7	���/�����t��MۃV����r��9SSӘT.W�&U��֟�P�E�x���A�@�_u��^��=�r`�X�w}����ja
y?����H���4w�
�����LN��1��.����V�i��;���<�Ŧ��to�j�p-�a�o���6��.G�**�󮰍s�M����#�UI �,n@^�I�?��w	Im.Ξ�����^h��s��yt���)}Y��=9����@řEchC���ϟ ��]M�[��<����B�j`�P=m�EDMI�|`5�.U�݌�茔�cRpJ�wb����������R�B�2�ϾK���ͩ�O����K�}��euߖ�^g��#�j��%m�Fu*��1����p�1,mpq Oj\��i�n���	s� *y ˸C{W�H�Է$*�Y�ԍ�m�bO����IqXˮ�Ϭ���ތ�7.G��	RJ0���q���VS_0���B�� ��y����yU�d)/.�@D�*3�/���f8��I4���[z)����Vh��u�Q�	������� �f����J��"Ħ �q�$��'i�,*Vz�׫P�MM�LR���"�*�I0�S>�!W������3��G�����U_�\���߀����Շ���~"x�a�H!!5I�>��+͚�ཬ��L-Ty����܅nL6&@��w�-���Q�*�[�oŽ�=�"^k==�uc����������u���.y�ո��0���ZHl7�t�B�"ܺ�5�Qof]�l���?B�>�$E�1SS���ڼ�C��3�U� �1 u�8l��_X����ޕa����83����y[<ZC���'XԳ����/eǠ�@A��B����ݵ�k�ƅ8�W��I��#]��Tp��F�<���7n0�p*�&B�y����j��H�\���v�J5m�p���V`��)s���=e�^="r��b�4�j����"q.a �,� �[��f�.ǫ��گc,��@';��8�hE`�9e��d�����xޥs�7ΈR��0��
�
��3T�_��D�:�:Nϖ�F���xib�1�S�t(�G��VPX���7�:���},j��T2��SyF��Vk���M�u��[��GD�wQ�����xw�U��I
5�S���&ӝ������57'^���?�[��bx9Cfc`)4���O�L��DM�/~?�v�jp��Z���_]��&S��,C�e�Y���4ñ�=���'y>��۽�zͤ�I����0���ܖ��h<&�됌h�*�V�S���w�<�
�O�n2fQ��+�<ehPD-��a1��Z�l��@+�0]K�w�D�g�_A-�bX�\BcU���P$t��ڳv3�Y��,u[{$���U��/GҠ�g���^��V�c@�B�ޒ
X*d`���p�/I-Ο�\%53��^�&�stǰ���V�;���T�F8MS��ُ}��S��M���x���D^��*#�q�˶�}џ_q�K~P�u�E�`���¶gN���mVh���/[��#a��LK�*^�eE�yU�f��@��fz�g�2�|�m
Vx�Sy!�I���s���e���jkc�,��#_n�s�}�L�P�mY�ϰ�`i�aXY����<�@͙��ڢ���Z�Zp�}��8z�D>�m���煃w-�0)���z����T0�2I��h�CL�Z�Ռ��g8��"�6�{W�>���2���]k���a�W{U�8-��A/^���k�����zg��>��)p��qD�ϼ��&u忲�~���J�M����� ��IP�	�tC1��{�]3ơrB���7U�!���f��	4�BwZ=C$�w׼�i�����������U-huS/�S<k@�"9���g�`�-�ݜ0�k�|	���ed�͠�`f�(�o);��?�y7��7A�KLr�G�	���*L�j���f´�T3�����A�~Q�0�� �{y�����9Y\|ǎ��Up��GX�˖,���(�2�]���ٕ�/r(^�����4�ADd�V8a�i����L�x��W�3���	=Q�`�'�%�K�x��SM����o�%�k��2s)��l���b������P��z�bU����vCJ<����@�Ò�l��$��x�"�0�n�ҜµSls�O���V�G�a�iP	�8ѤXY�Ƚ���=4k����r[6ӣ�C�BYv5_��n�4!��蒛�h4�����9�g,����6�`���"��0)������Alz�|���v������J 	"Yz�^�����X�J�3c,օ =�����9?�]�	n8�Y�6�7v���rr�{<3m���a�1�e����t�㧣�hl��r������A���lWv�D�@ex�=a�^g
���ݙ_�N]T+�I ��'�����>�"E��I�8��z�4J0s*�n-~�L�s	KX�p"W3�"��~�^��X����q�2/�Mj�bMS�� $��bY�{�^����'��i�@K�ܲƓcu�&(K9�1�`)��\(�,�'�R�}m\�|���O�_��^���=q�d��k&o�V������Ak����w�º�C����7<���è�uG�71R��<�Y���*�x��j�p�2W%���3�<����x���	8o̍zH��l�g�<�?�Ȝ�5xp(7��U%>m�)�_j�LR��%(e m&�5��2����e�)R��$���0����$��l�l9�<�̯�#��~W�NޡU����C���;��%��؋r]�
;����a�{k��4�aС8\��Ω���_%Rj��k�6l���� p���"���)[av1�軝�z�3R��ҘR�t���ƚ�����)�]'����NE(�E��g�,�n�^���ly�T=��dPf����i�ʆh*Y/_�]c]/��φIaJ���^۩Y�dG�-a~�lD�^�G�k�n@F~��(2���)Bϛmi58���#�럭6 Xmϼ	�T؉�Zݨ�bi-m����jx��+��0�te<�Է>'l I(���u�����HET��rE�@�&����{E�ᒔ�}J�ř�	b��U��\U6�)f	nn���w7�IO˹�V%=���>�\P�"?c��j.���u6s��|d{Sv����!m�T⋙g��XUl��Y�if�b�B�NBE��Z"�Y��� //���&��Vݦ� �w���޺� ��#J����W��U�j��'XH�''�?��o���c��C��2�� �8�	,�+���hךS<�Y6" ��:�i����o�:=�y������|d�/<�>r+�ApE�
�q$��V��'f�E�!*Dx�{���g���i@Rj�Q���Iy�.���Dā0µ�r�]�.*2:j.�gP)Vd
�t�43~	�L��*�?fp�_M��4��Y�x��
�!��ټ9���W�D$Fs�c��Zi׌����fMa�h��vŰ��j�I]g�!��W�7l��q��ԒK�Z�Z |��K�����_�+��[E~���[a]���4{��lv�lx��=�G"����"Mh$�����#S�W��d��̽�F������z���妞0�;� 9zY��{i�m(��Tu3�7AH��D�F��AQ>F�m���:�7LE­�G��d�բ��Ù�}�[|2�_^ C�͌�S8AD��n�v��'�6t� ��;���~���4��a��?�w�s��$�@^���"؀c�����p�_�f ��W����`Ud`��������qu1����>��9��C��C������c��)��ڹ�",���O�( P5GR�nd�6�Z1�^÷~^*�h�7zX-ojSȞ��m�_,���-�����Y˞�uL��9�M���.�q�}�/��HU����PG��9�u���b�޽ӟ��j�F^�T���V�����S�$�jy<���H��}=�Ȓ�4}b��}(����X��u@{m�|��I��]�T�l�_�eL��C��B�A28&�lK�C�_�UG.��R���t�W�4�'�5<J�l�ߧ�Ͼs�3�ryg�X�]-�2x�xˤ�X[3�{6��*6np<ԗ�ٌk�nT�<u�P#wp�����jq ,�Fu�H�����{��A0�OY�0�z�k���H4�yZ�!H9�h��M��J�A�ޘ������
��w��=%� ����S��vj� w���<�������^��n�ȣ��_=W���Bu8]
*�^´�c��(D��K"F3X�>����Mp��׼�=n�y�lD��iT�i��tđJJ����!\�w/e�^�9�+
S�_�DCz�BX �d��F.�HD��k�=gC���4�>�+�������RD�S���*����R�>�ّK-���)�V�(vixJ8���vۛ�u{����������D�W�ƨ�f�P�]Fb�Б�3x�kv ��!}'�~=#j��p� ���#�"�%����0�P��`��&���?�2�b*��@��4`��Sfpf#%�f j�^�"�х��o��߼.<�� *t,�A}�� �e!�7�JU��AW�!ޣ2�S��NJFM��)^��h�<Hn�[�'�e��S#�w�:�����#�[%����P��<�b� {��ؚZ,8����%5��� �'=$�H��΀�>��[�܋�_�vqu�؄�fa>��yPNWS%��JZ�]��������QN��oK�A@W������	�ӣ`�yW��z����(ЩN��n��N q}�>�F��Ź�7�p��A5�)����_��d�e��R�S�>��ŦТ�b�H�K��l�8A[�v���E��I��T�Ł|z:��־�S�2!��6VP�ϖHd�� Xj�׳�s���2K�lP���ѕ�������E��U�>���3�]��`�o	�`�2�6cq��վm�i�+s�xz��5��h��<��� ��N��N��$��4��1D@�!U,XW�0�=����l�����y��X\��X��F����,m:	�٘���&&#�@�Ś�!����|�{�h�~�Ԩ���C��Q�L9	oV6�tm[�7f L��)���8����;3{�}/B!�N�I���w3�uu�/��-�L��p�P=}y4�p�p�_��p6��ŞT���ujW��d�aO�&�9X��jd,k�&�&� �٤6��NA^~y�j7jXZ���U[�WE�;��HY}I�g������Ă�y{�1��}B�^#����8�&M"N�#���DB�|ƾ!�����dd=�،l|>���q���1��~�~����b �Jn�S�+�f�um���+���[?��`]��0^o��"	��l�U<�#;��b��i�1��r��j!y�~2���z�����s��<ȴ9m^Qq�CJK��p�!�.G A9BH ��@�������Uᝣ�ٌ&+��8)��i.zKV�MOp�Z��%,��B��d9�����p��{vp _��j�����N�.
Y���Xy0CX�R^p����@�y]Z����cM�K��1�k
O.!�5
)s߅��4�R� V0���-�;��}z��'��zt[�?P�f���-�v�4�I�b;��夡J6���֛��@�챊c��]WV���Nֶ�Au�����zX-��p�X�2U#���w�-{Dg�N�)��iH_��Nd�ޱ7|ɮ�i���e3�J>˸��D_��es%�l
�R� i�m&� �TMQ�׵IDڃX�P��u2���ř w	W�Yu��*b	I�B�^�t ��퉀e+y+�:��A"�HVl�]H�-舜4j�ʹ�F%��6w���!�a޹��ힿ���Z�P�]=��E;ܹ=�,a�7�6?�p�缰k�W�H�ΐ���yWf^ݱ��-FϺw���ڢ��E�k^�M��k�i��2f�T�a�����h�W��5oȪ4[��ʀ��8(�1�O��+��`O����I��v�	k����J����vސ�Yɂ'^��;�z�W�%PO7�W����:�̠�-K�5�r����jBi\Z���v%1+�%|7~LD�ttO�g%"���{��b��(r�O�<���L��;��c����'z�Fz�t�!��EXR�g���9�G���X�U�#��
��i�Y �k������f���l�����+���~,�_��󙦧g�a�#���LZv�hIa��0O�[���&�ue�!�L�4���@���˝�b_�+�ild��?���%�zo'���;��YS����Ї��XI\@���������#�RW�4Q�������")4[j�.�Uo#%���O] �U��ۜ9�m�+�rE�{��b�:d�w�y7���Ĳ��l^�������a&"�4rѥ���Fp{W�z E��A���%�q�\7}�����,�X�Je��1��4G�8���g\��i ����U�Jc�Zf��E(���;�O��D��-��|�ݐdI'���:������k^	%�%���[Q!��Y����B�0���]�,�q*+����zC4�tQE�����%y�2=�:�#�}[�,9����%
�P�F^�@���N�M?,&�G-����-�lGWB����X8�_���>�t���/���gpJ=���T�2�_N��@�S��p�2�ދ��W�Zr�cb'���QB�a��t'-��h��}��*+x`�и��^?\cn��ğ�@���Z̫��<�h ��v���+W�}�ެ4>�*��sk
���\	U�aq���R�q
:7�lC��*��<�_D`��c YئZ%���O¯���6<G%�u�nJF*���Ƽ����M��M�WLY�y�|��gmeX�url3;��^)�\�\�64���M)x<~�?��w���^}+�4�o*�����#��!
]VU�tU�FF� ��u9�F�l�XN�^��F8�>O�!��L;HP�1��Aqb���a!�h��#?���AJ���fi�5�"r;f"���z��ˏ�� q|��abЌT>��/^t�-��#
�c�һ����2����3-u[���Q�16� .�����P���K("R�d:��[w���Ϻ���D��7M=Va;GH9 ���|UZUy�/�R�˟'������`�[�������kݩ\#��*�i��A�����6H�DY�F���*���BdD�DD�F�4��;p���+j�X�-b�-�V��aJ/,C/�%��L9�����L�_�akR��113���Ё�~)yt���H��jY6C��1��`T�B��N4��Y�VF ����2oi�w�P�C��2�1��lQ)��ha�	h�Q��OE����F�i[�A�����i������xU�vvw�\���v����P���*��X��o����DpyS��9��$�����]�+e�������jI{��#�nz_�1��I�����#�)zo�&���d݃�`�iL�c��?.��oj�69��e����[q-2;>WU��ŲX�=��;gq�M}RڀOOj�&���H������x�m9�I0PU���$,�%�o����r��|x4u�^bB�3�+p#��YF-4��6��6O3�P6�mL�6��ieۑY��l*Dw���إ��n.ʃn�����x��_�,4�ʗR�4$��=~�:"{�k��x�T��@[(<��vj-�)��ؓT�� 0!�+�­��j��K�+i��3&$f�X/�le��o�������fu��쿝�;U�灳h&���><Ud.%�q]+�n��SS:�u�5jZ)"�H��9 ��;���@���6�`iSj���̐:�ы����=�|d�I1�k�6��S��B?c���e&�C����zͰ�@�'��"��@��<�����K��4��y<�3XK�vsS����b��}�ڤ�OG\���%v��Tk� $glem����X�Jbb�����^x� "���U�FΦ��=	�<{RY�׺��\�N�>�:��`[C��/r:#���>���K��s�xU��%�Ճ'x�!�*bJ)��2��r�u�e�-R�a�%�Z�b��0:�pK�&T�X#l�O�	��d��eb�4x����R��4#�+��v�<�ϯ�T�I���iC����4)�+��&���+�+еm���C��hB���T�-�}v�m�,�w�KQ�J���F|1���]��^�'����󨒼e΢e�`���X�*#�ר͙sܨOFP��f�����.���#g�!rۂ�ā,�\b<&iܚ8�kź%��G��q�n6����5y� *ys7ö�]�{V`/�_���`���s�G�r��C���Vû�;�2��X=������?�F���qIq	�	�5�+-H�[�<H�Y���k�@��J��3��=C:����fs�_H��G/�Úm��+D�A��^��
`�������L{op)��<��J֣HK�8!!}]Q&KX��Qˣ�?I/�aA�<�$���<�#��O6�)�Q A� ��#~���O0{Dd�Y�*[��������>e�h��[�k��+�&6~��6`&'��(>q,R��P��m9��A(���ۧdvº���K(l�g���Y�ο�Sb�W2��J6�Io����M[�����hЌ�lu�~_�|�*�|=z��iJ�O'���qb��?�Jg�7�ۜu�?�bQ`�tym|<��j��=��f�T�$yo}���w2QԮ�?ַ�ź�N��s��������t��O����q�3�7_�Bi�ߨ� �}_����F�����0��.,�`Ǆx$/J\y��Y(o{�~9��@��F5�N�[��cd�Q��^5U�D?+J(�����bQ���J�zA��<lw"�S��m��)�Έas�pJ�lv�5�=/׷�s�]�S��b�`?r�/(	�������H1�����b�#m�T�I��x����0~��z}؀�X��|X����Iu���9I����Q�j�b�k��mj����k�c�Ae%3ˆ(t&Ǖ�5~�qjf�ěVA�{�i�#�U�[Y����)-��u�k���.>��pFbV�k�5�`5�Y�?�ą�xS��o��G�"2
��$����0�D�y�a�v���될�l)�%
"4)ѯ]�B��-@�[��^�j��6/�'"�(/�n�W~��s��LbH2	�pQ͍�I׏~А3�,ͫ큕���.��M�� �$�kV#�dK��5�i��~�VRa�	�9v�Yڱ6�,��K�Yل�YN�)��͸f����� ���@��js�&A�)�L�����ٷ�f6/��<0��?�\��f��(I�l�	+��^�jE�>�l~�eX:��D����?;!��8{_=-��Sڄ+��̂�u�����\�n��d�1�bcF��0�T��pD�� oK���/ꆊ�~�&�$5�.�>�Hy��W.�@���튟���4�<�_�8E�=z�����|��s$F�y�x��o�w:� O#����Ja����F�2'�S�sZk�R�����IV�N����*d%��5a��7'rf�Rvѻ��E��2�5�lk6�[�±&�R���a.SYC�$Lz�����C~@[Q:?T�)�x�4m�ɤ��?���Ü��#Vp���.�[Bp�檬ds�&�L�z���Ϸ�|�b@��B�1G&�t�o�q$�R�I>a�85��
)d?����rZ�W0H���Y��;����a�=�ǾU�JȠ4�ջ�DX����[ؗ���|�����2Uaɘ*��y�5쨸�_��+�u�C���w�J�AUJfd�"�ov�x�0Q�J�T�@Kp*�Ԫ4ŅF��({{��g�IŇ���H'���iJ7��̌#���m1X4�D�u�ЖL���>GΠc<F/�W\	�u�K϶o�[���MTd�^��b:�}��i���w��ir��Pķu�>G��N�-1#��w�R`��|�O�xP��N�o�(��Ib�ډ��.��*֕�ˏ�&�����J�N����tO�n7i}����oS��F�&^�}Fҍ��]�	f�؈<K� �6m����@L�끛��m-�H��L�K7�K`qA������d�
Nl�����l���1b}�߆��C
}�?�.����\<��,�@U'g���W�IL�-��p�ZDa�K�_@��Ji�҉��H�{���"o��Ѐ��@th����d��R�&đz]*Y��;��<���m�%��
�:����5���>�&_2N�������^�ߵ߃`/��Ԥ9�F���D�R&\Mc�w}��],G߀:�C@��=�Q�4���P�	�3϶��g1��[�Q�khUcR�5b�|z�rQ�%f�:�ӹ-E����u�L7��bu�{K��_��_�����@�1.{
��
��XMڻ�@�Cov� ;	HDc����L/[A��)^M��J���W��-�5=�YnJwj���퓏�"Q>zL�Ӱ�SQW5�������H��5/Bl��j���-������߉r$U\��O�����K8Y���0�R%����D/�*�T�a��J��B��,r3aQG�n��ݴ�Q�D�H�P�e����`$�zv� 7 1P�I�i���2ĵq|;t�}�/[L�1}�f�Ț[!�Q��u�#���������jr�o	Y���o��h�Au������&��v�������c{qM�"J���n���6���Ą e�г����Ld@�M0`�R����!��r���p�@��J���Ev@؊tߟ�ب^�͂J��~д����TU('�م)459֓�f��>��w��n����)ZL�F*깾�YZ��E�
Hq��1���J��BS�����a饸��a@o�:���;c�4�|Oǟ�f����~6��{0h�B�+�5������/�WШ4�"LמMiY&,F��	����V��Ë�+Hq|����2t"{Ƒ��Z���'�h���aS������%\<&ӕt����)���^3A��M���B���y;�Fg��;�6��������ԩ"��'7Q��iy��	Zh�¥��P����K�~�k�!���b��
h���y�H<����(Ο��M6�:o���"$�C\���`w��P��Ȃ}���Pg��{��AYJ�Ͼ�o��	e �	���U&���6Ƞ4(�����
�y�����.�?���u�`��[Φ�h z��57��%���n��
$�b8�[��G���c�K%�Yӎ���63��nV���t�������e��o�Ь4o-*֔����@��^Y�(��i����S�D`�}.�X��h�{c4����p���sí#�������3�3B/�Ɍ697����hZ���a��@���B���:i�'�t��R�x��3�hsAW��o�M��RW���1�p���F�7˽��r>��I�bw�zeT��B#�U����N�a���(l�s�cw�b^�F"��;
��'���9��כ��d�%�J�+�B�p�:��b��u��#͔C/���aT�X8�"g��n��T�B��o��o��4��3��{��!��h�!�5�m��iyiO��4�u4Wʂ9DM�U�b_���#̘s�^d�1�B�YnI��s�Q?sV:1�\�h2��$K!b���U��oA�f�BCb�6���]�Q$S���&�Ny0���=��?��r�faA=yl8�0Fs�"`��+���F_�hdY�$��7�c�����gw2�X�d)����L��²��Ϫ㊕L<���T�2�����NK��7�Ʒ��?B�/5P���s�����-�1�}�
�k!x~����Hc��k�Z�S|Y٥�~5'��jGΉ;�d�Ҋ�MLq�|��f�G�I���w�բAւ;3P�ÈM,×Sr��m@�ո�k��]���JyO���A����`��(�ǭ[�>>���ۙ�&�E�$�Od�2��*���|%���*|ME��^1�C�]�� /WT@�(WA�Y2���w��T#	0
̝��T8fv�H�+Ӿ��@�0��-�gӊ z��cs]���aC+����RF�9���ꃓ{�_;��N��ƒ%�����k�(!����E�D88����b�f��;��4����F�aܩ��i���_�Uұ��P��X���`��$
0|���:�
?D�B�9�|�C���C��-�����ʊX_Asf%ڜ#��ذ�Y�?��D:�1���w�F�d����[�x�w�p�'��U�Y*���[$%lX�kiQ_��AD����_�;/��Q�s��%;���틼��L��/�O)7�������镥��An�?��O��fnm��q���a����x΃n����=
�;��V'�t�9�<B�Ś�*��F�N��c���O��,$	f��{o�]8���h}b+�[�G����HF�L�ɷ���\��	Sp���%Q����!��	s�W��]����rx�0N��U�FpҌf�L�uk�&2�+4ox{���^c�4�1�Lb���/;���j��+<�v yٛ�$^��6Rw=7:/e��5
��_�AUJ�N��~���B�)?�{�x��:%�ۢM^���8U����Z�PKCS�A�=��rulwK�Í��꘭���9��~� ��պ�#��� }+W�g|�\ֽ<�,
1�8-���3|��>��w7.e��K���o˪�6�r�;��������_��� x=�V���c���ғ����~!�0��}A�Q��aN6	W�ٝfCO�~��$�5�c/�3��H�I�T�?��B��E�`7@4xo��t ��38yY�|���������6���-SU��p���|Y��
��G����+}��CJ�	��:ວg4D2''J�wJ��Ѥ�n �Ȼ�Dޜ�fԲ��<�uݺ=����C�k��'��z�gZ^�{��#�x�~�5��v4g���<��p���u�~��*8��41�x�R6�)�u�/����/Kip"f�����7�i��p�ѿP]5:��N��`a����L�06�D��C�!0u4 ���]G�@�-�)�<�Y�4#2�P_�o^DRj��ͺW�i�L|G�<8��&��"J(�f��)˅f��*�ҵ8�xl�ը���Zu�f-���nФ��f��M/���j�2�0D��������Z�#�����wc�]bULz�]����-�����d�k�_�im�}��i!�Z7f�t��M,B��u�`u��UER5&V���G���#U.��܉gd�+�|���l�i'����0���*)Si�43!�E�l&J�s��c쩐ӻ�+� ��0�f[t�+����I|=�T�b��k������J+��>�@'�s�����̎�Ih�iqVKo�Ɔ-A�>�C��TS� ��\V�MY�M�e��`�i�4s� \�ܪ��0��c����Ũ��w5����3��5�uf�k.3J~���N!�"^�ס^�qu)M�S7<�L,������|ȷ�ۤ*�V�)gT��g ���c�EE� �HY�7�`����&H�M��V6�v��YF��u_��`�"�������#<.�܅:D
�l7�9�^�;�����1_�k�-q�bM�f���#�HM�)z����eG�+�|o��SCu]���� 0&[Li b=�'��j����sD)��g��^�]��1R��A�Q��-�-�M�5D� Qao�ut\�(�H��t?���2��h,��
 �=0���(~���01��r=z��n+,s<����18a�,�4����I�'��:����p��Zj���WǮ�(bH��n�yA�,�0C|�z��=$��N��'�#���v�c����V��j�dq@Q���fG���)NNx����Eo)�EC�&'�m���]��EC�U~�����鳿�>s���l#ywCWD�����V���@�6Xj؄�5H�k!;WtL�B_ ��U��2��S?�G�Ilɾ.�(�rZ�O>����d|�g��t	QE�^���ta8^�wN$еrF	�0N��WЃ��՟�g%Տ�b.m���N6�:�sUOE�k��b�q�s�C����)���Ma�3��݊Z��\G�{{nc)���6��hg��`H��~�|�_F�7�	�q#�vK.ٽjj��H>��iw���6�N�B*����BW�����n_��̿ᚦ;DQ�ٔ�J/ʇ�t��m�?{!��98y��1E�w�}��uR�}��1u��M�I�'?$�.�H:8�0��ʧ��*RA=F��=���:>XDGd��~�1�Ǉ�	'����L\�g&HTak��3^%�$[��8�^��T�H~�!Z���Т����Ëtq�8���K+\z_N����]�i�C^�W���V����F��p���T�y}?"_���M�r��zN}F
$j���ߣ��$3��+,X��M�#�j�8v 4W%7�,<
$r*�� �r�t�7^b�Zku���#�~dA#��3d9��La�7U��}m���'��i����snrQ�B���`��zDmg�ܠ���eB/G�.�S�a�u�δG�;���ɏL��6���x��g\]�^��΋�E^����#����Ɛ� Μ-�rȏ�饛WA�ac.���{�������-}$zg�s'ꥡ4�~K��B@�^���*�A�-�^>ɽ���ʨ/�[@\��0��GD#�R�A�˷'��=�q ��ԁi���W�n	l�q�G��p���0��������3����H�c�B�50L�C�(�m�
#�w��t�ҷ�e��ߑ*���=�����|�N7 �O�%#Fu�SU��Q&�>j��g����>��?Ŏ���$����<��J�, a,r���������&�l���ӧ�+��� fi:~��+-�!����D�;�V�S'�PH­��\Jb��}���@O5�p,$ ��]"�
��L&�r����(�H��z3�A���?u!���欣��L�,�$�/:*�R6^�0S�w�J$=�`���.����o;�#�^U�`pk�ګ0CK�t+�-�#0�~2i6{���s��%[�jZ�)�넛�r�Zca�� zK�&�1��KU����8�/W]������|)1�ek��C2z^�a�<ڲ�
J��s&���7g@�_�����śA�|ډ.Z:������]ec �=ܜs�<TZ�_��#^����5��q�ye�SD��3��U�P�x8���h����b�9��1~����7�?\�����t�7���e���Mt���O�v�]~�W�0Cy�5V����r�naE��~Y��T����9�Y{�ݚ����|9:��U�B-��_۪�ޯ��v����V�{�?4��KB��u$R����Y�ش�5DPآ��"�^ ]O�.��Q�1�ܚ�+z!r�i?���h50�F�.T�z��{�c��(�J����f��n��G�Kb��HUh}\��˩�{��������a�3/��`b�: �\X� �ή�N��%kU���?>4�Y�ܩ���	E��.�0Gk�oM���(�����ՙVy�����N�R��: --����g�%f)$�k�8�Nm}��J���t���^߯��y��L̤�%x0��*���
x�	m?���E�bzu���U��lb�ƽ]h;��
�@>�C;eqV� ����rU���xC��ϑ�v��(-�;�r���?���/��\J;�4�C��;��K����"C�p��(���2��+
��3�5[��΅�=Β�����B��0
uW��d�'*�ty2Pj1
i[�#>����(?�yY(b'|��q��ŉ�̀�,�Ҹ}��Ư(w��)#�6�Y�lo
ߧ�2���"yS����X4��kѫ/��F�nZ	�����W�y�m���<�6��� y�7v&10�XͥYa3��v�<F @j�'g�3?�^��7@O��
B�b@�ix�ҵ�������+�$���޹(W��?k3�������@?BlU'�CT�j���m>���<�T��K���.n�wJ���#�;�?����ìƂHY�z��!ъ�q�gc��b8�y[��r�ɡ� ��������x���m�$��U�]����jf;ną�P�FP�]��������\!�sL4�� 8����,<*�x-#�����-yۛ
;�=����4����zvA}�Y�(�V⍤�s�]2a�4N!?���H��x�p<Ms�e��m�_y�@F��HB�o�37�O��Q�B&��fc��CSU���!t�0����k�t݇���N	W��_p�;�Hp)��?JL^��)����e���;���K�n��r��W�g{b\��)�*�<p��E�7ǝ�P͆�X��x`y8m2��;gp9��s�3@	ޑ��I(���UqG�2Yo��ro�9�B����� �*�ȉ�<��Π�`��)!��]aX�[>���GX����Q!*¤���z�ߦ'_ErmF&��>��玠%mph�)�u|Xg��j�w��7'G�Z��vz�?�=�V� �y�B&%qR�3m�3��҆���Y7�7�s�^�:cE��c�%�6��cČ����KZ�8����.� 󫜝5�v~8f�^p$�����c�d5�n��M~�N�����P�����0�8���O�5J�\!��A�o(��-ϳW��`����i�z��1�q)Z� �����h ���T�����C�5zv��������?d��� ��æ/�����}?;�/����$T���˳+
B[K/s�3OS���T���,�ږ/5�E��OM� 2�'�1� D	�w�@����)���L�9B]<�n�oh�ˏQR�,TCu6	�C_���Mǽ���Τ1p�~��{0Ќ�Ʉ'��p���X��a!�$g���zS��5=ivÞڮ��jpC����J�uI�0�N��zP\�ɷIYe��EO�������(&3��[j^j�!��t �Xϗ� �[���d�bq2����Y n
��g��a4@dd�O���|T��!���=��P���]Tƞ^P�f1�I���Hվ5Z�ϗcW�z�~���z��s���ʎ�ij�p��˓�N�%��x����V�O�%�$WփYB�;��cIЦ�'�I�j24�E��`.�J�ɧL3�j/������Ф��aS����2�`������-��9Oĕ�����o�5��+%Վ�G��h�0&$�OP�nnK}]w'q�i؀B+�A����1w�q1�TX˨�$������勂�rG~BOՌ�$���f��j�)>�ՊF��a�P V��y��s͢�K����M���)&��_�b`W����J����^{�,Y 59oŭc �c2�����%�oPĳ���߇��:�K��j�ŗ�.�L�����},����-.�:���Н,<��c���i+,v�XHo"���4�	������@�������n�s	�f���30[�t��ky=�R7��htؓj�U6��Ej�=G�"��[���=����ڦ+q����}��y������g�Jn9+ɚd��c��	��!����`�E`���s8ƫ�J���z>$���]�4�Ԭ�",:�sz�vKJ��* ����,%f"�Ͼ���c����U#���3�Ύ�y�'��G�F����l�c`[���吉�c&Q�_�W@� �+Q�>uΦ2ږ�ڨ1�o~�}�F��M�}P(C�~hS��{�؁ގ�=K�������^qy$/��bԺLo����2�Uu�B���,���bHﲟsd����kZR3��V�����լDq���bd�ή'�5l,.b�(�����{Mw��f�$&O6�r�P�2<��R��8�^����'2�oq;n�'^KC9��O4�
�ϟ����ʘ2�)凞pE���V\���/���l���P��T��}��WU�4��;(��zIa���|iK�Jس:s��7;
~�J*nb㧾s�H����#�E�xȎ��H��!U���kB�ww�!&%D�}�1��g����z� N�6w�=�#	 WJ
��Ϟ@zFZ�p��d��g�力�5H�!�&/4����r���k03��e�{�8]� �qf��nM�Ya � &{�y�:�L���͞�={���������ӊ�2d^�yN�DC��wR"�Қ��뢂��$nA��*��!T�/9j&$�Z7i��y�qs#젏7 QGhh���V��qC�v
��إ��o����;rT���x�����o��k!V��-�l���lVϣ1wZwi��F}AϮ^#+%=��_Ř���ހdZ��u�#���e]T]D���U��,��e|�}1&y��Y�xO�Cg|K��$���>���P�i�df�$�jsCvȏB`��]�£o[1��M��U+ϳF�K��0s�5a-��o4��/W#�d��w���e��1>�%�qy�zuq�=J�(Y��lHvQ�Y�w��/��zo�+������\���Lٲ�~^��s@��`4|���e`�}�Nٚt��ʙt���li>GΦ~T�AyOC�r���}��o��R{IA�Hr[��ٴBԭ��]A�gV��e����x}�#B׸��u�P�S'p	�ٓ�S�C_G�w��ͷ���mV����}��j�!�/Ų�ҟ���e���G�B�NE����_N��1cl7���f���NŴ�}�䬶p�KFJ4� }���@�0 d>U,E�
%��hv�E�M���1cY�%r��_��:l>�uur}�̈j�5�޸�|�b\���ȗ�`� =gr�k��eV��#Ț���?
�A;�ב�S\�J�v����#7�	&~a�p�*��� �ƽ"���u=���=�sF9�)��m!֔'��ЛTdFm\G({Bz�˩�龪�}h�t;�%b
�cA9e/ń�f�$�ю�����tJRA���hM���D���N�����q��ɛ�V�Ȧ��{6�&w!X@��s�a�L�_�&����wE�-�Z"�p�
�~����^��9'W�1ص�(�o*��i�}��E�.�@0���>�|���{@��#�Y>� =Z��S_�ݹ�J��/+v�����]�ڋ��$QΤ��1$�D ��fÌ�cG�T'�y2���i�>�����T=[E1@�9�%v_��Y���{�6BkV?���{�r�I�un�5(��<0��JNמՔ�X�bg�,ϑiY��t�@�W�H=�[��{�٥]��.+<��8D��H��5LI�l��i�btG!6�(��afN��	waN�Z�t�Q��HP�~�DG�z�S1n��7����G��>[��j�����D�.�&���G|K�ڈ=h��,����у��9�f������&��Kk���@�5t��B!Q5���X!_�2�!e��;�P:o0d�Ϊ�r�۫�Od;1���Z���l\�3>�]��B@	
���c�LY�߭nl�o��~|�-�O�����4e�}�T\B�_���n������c��{��oU�1��:}��4��À��-�y�،��h>�����i�����SzTY�C�ꃜ���	�s~��l+�D�N�x��پ�x?�뾝��;�������\�b�a�Rf��Q	���Q%��(ee���ʠ�!c��K�e�?���i,w��ȦG��l,�uK����K8Ä\T�.��$d��O�n�q,�T��~3w�p�K&�+O]� �3΀�G[2�sR7�<�����)c�Ze�H�,F���DW ��C!b��x���N���(�� l��!�K�Tv?���j8 *�G�]d44��c��g9�ب����}?�m3���b�4��#�),������q�� q�'a���/8�UR#>	�T�[�S2���f"��c�U��@�<|]�'[������{=�<9��)�)'K�� ;yz�m��x�MIu�ʪ_��I�Q�>.�x�J�D��M�K/�Oօ{��$o2���O�od`��2�Z�3��׻�Z�3�G	3��MM{fL-)��d�f
)����=�:�/"͇���>�>>]��p*E��y���P@R�m	!��1�=�0��w����?.�[}�5rңVd��9��n���gZl=�51c�b��e!��jD.�����@(��UXO�c��a�&O�ƹ��zꝆ��2Y��!�D�@4���5��>x�D�L��z볚�I}�����3���[I�pp�wO��|,�8�N�0v	�z�a���s�����C{`6������Xno�ճ	á>�f�݈5s�c��GiB��+�ih���x�d����J���.���V�o��+}+�} ��}�i�H�0�ne�zǴDPҥ~��ˀ, zh�`��#���P�zZ~7,�$�x \�� �-������ٷ�ch@�s&��M��_s3��Y���}]q��?&U�Ǘ�0ٵ�GWb�����zm��o'.��7(9�P|f��&)2�gr�~2w��/�(KK�7��]�I���ఫI�������(��Y�F��)���f����y�K����������Z!��c�~��54ý��]��[�����A-�P���M��!�����GѢ����1�.{ҩ�kn���_W����G�Y �^��iz`��'������cv]�~- ��<xd8�M0ng`8� H�\��*�$jn������ɡj����'���i 
(-�d�k�j(��0��EA$&X��IB���O�;�J����Q�]�����PK��շfE����Wq�`����Qz�K?a�_�?g=���D���8�������	&.J�����'�E�e+d�S���{��Yc�Bьp��G�J�5d���܌����s��'�GZ��J����c�`�.lx�l: TR׻ �-���9\��b�f��I�� ���_�	hZü����8pk��n?��*���s)F�*�q�p�ѵ��&,X0�v��?�PF��s�����F�a�<^cM�"&��J3�|b~E�xF�<0�X�U'ʙ���Y���Q����i��;n57���nGC�^�5�Z��q�� �3�壹�n����d�8�;]��V�rr最�p\ �hR�c���$���@.'����(�i��rzx`H-:�T�]B7!�'�xK�
*��<'xHuy�{�^��+P$��^yY�4?٘՛a���A�Mg5^�Y7�'��3Տ��r*�	��ڢyȭȐ�����qi��+�M��n��߳.���S��*�}�^��pq ���&1f�Yl���#��*�9���9ҍ��
ĝ��l��I�~Ѷ0-Ѭ`��b�s)���D&������0���fV\�Y`���qܖ��2`�]�'�`|�\�+�V�$���^^V!A�]�1k�n�����R^2�@G�{U��MIj�u�W���DiyrRU�5q3����]31M�9��MV������Q~!J��H�!�Ȭ�3T��B���T0�g*� ^���|�=N�/y��M�,�IڊB`�9c��Q1 ��>�eK�R�z.jo��r��:ws,M��'+��4�+��n g����� ��l���8����km���l����(S�J��l�#G2=�a��(Ǥ�!Ұ4�BV�K܀Ø�L�j�F�)*<&��ȓ��)]�X��n_yKi�x��,�_���PӋƙ>q��=�����*S��Z�~=IK�D�䰺��<���B_D�e*��P��hɿ�(���>f$����em�=������|)O��ǿ]�x��|�/��] ^�=4����ޮ�����Y���.�m�������p��0��_#f�*N�`���0_�1s3l�I�J36Ǖ�2�p^�fPr'��Q5L�:F�����O����f����	f���(�`�٪:�5���}�'��n�曁�� �@��j1+�4�<�CVK���������8����BpGцg1`��+��G_7��
�\WQ=����o&qO?}�$�z����3��^j�p��#�d��W�J��� t���~#�ATd�L����,k���(�V[�_�z9b�N�<@�����n��ag�+� ��S#���n�
�v���V����d�,s	�NUH*& �+qc8�
�~��󈰕Ҹ�"��v��1��K�t�}����ހ���$��#��/��BHi+�aS�UV��9�p;/��\�Rg[70Uo�e�p��+'$u\T��x�e��^O�����v\9��mZ�((8�r�M��L�``5���B�������lj���v$]�YǛ�{�?�U+�����6����@���s�=��G��H6{��b�ly�G杦#�d.����EÎ{l�q�R�-��W�)o�([Ԑ����8�F�R{sW]H�*w��c��F��;���h�;�i��[˧�XQ��2J��-L��������� ��V_c�j�^u��|6q��/��T�3��V�mhB��dsAHތ����m�����l�ƚ=��Z�_�u2V�f��f�����SQ�����M�����$"��]��rC,r?���`)L�1�sp�E_ʝ�t`�����ub'`x����"o��bn��s���~XA�9�0�/���j�`��%f���V���@�a�y�%����?�� j�|�.@cO��W���G��d�>j���H���հ�����$�ёp{�)�֥\÷:b����(�j��Cy��,���*�	�j�֋����Q���a��$��>����b��)��vPw���m�����E�X�pl����:ҠgDA����������+��c�3�
������ϖ״�%���/]>�ڳ��#������n�X��uz�fe�9X���'��;���7E�{��̊�����W[��v�Fٗ�x��V��,9el�Kx)�{�tO�9�
����d��؍O�����]ə���������LP�%�,��<���>�b\P�:���u����Q�, ����Պ���o�G/b2��D�jGLLRUj�J�]1�T����>��qi@}���ج�)X.P��xl�.<�#�(���$e�`�D� ��}��8�<���eV_�z�:�w����=<�	�0����(Y�H7:����6ʕ��5;`ܩ{���(�4'd\���j�-��i[jP�8�*+ʳ-L ,&A�ra C`3i4q����-0>���C*9E�Ru��-0���7v7D;���Z���m�����V�Al��^&y�d>?����l��J>����?�u���&��^���� 3B���2�����9!c+E6X}���W� ��
������⪄R4��!=�7C����v�lٟ/��5EWz���}d� �ۤ43��9Q��g?��#N߰��萢����݀D'��}U�"V{����d�zWR6L�B,�#k��M��7�|AouE���>�=�k�vd�V�3�{�-��\�U(F��
y"��@��쵮׺�4h�Ȭ��^q]��bFq�u��W�)[0�4�ޔz�+�6t&<�~LA�v��n��PHM��Ү��?gQ�[��t���F��HA°��S9�ß�%~�nj�ڥ-�	V�����9�<o��[��J�@��u��e��11�����Um6�ˌ6�̔n�Q�������ı��r����e/���&������h���O�p2�4>t%Դ���pV��ZflҴ���{�0�>/���\���،��X�2�WΝ�sqv�\����J���3�-=rs����V�J9W9L�Q�u;��	T?m��; , 	+.�T�+"��eu�w�6B{�H��	�|��ZOk4W�+�3���2��u�^T��g
�9	ˬ!DYr3�r�򌿞b��aS�"�����6�����ɪÉ�[�$v��h[�WM.(�(�E�9��po��������as#'�?@�8� ×$9,Ne���:B���ٻ���9x�i��� WXWgM���ƸeMD�_u��4c<W����$�n����t9!�sބS7����4z��Xǰ�̤�c��iFF�7(�F'�9�v��z�� 2>�z�c�EĹ�,�Q+1M¢pCU2'��={oh*H���!��؇���NDF����mV�^3� �5�ŋԷȏx1d��T���A W�����ĄS]��Vb��f,Lu���dNq<��ϋ��݀IF��ۤ�,q%I���}�I�P�Q��~P��V	��g>?�/I����	F�&�v��[�s����&*�nj��E]�>9�W��}�g/�.�_�6�Y�1}��>o>#������Cq4d>ťd�W�rD�%�d�KYG���$+0��2c�FS��h}c�q��QY�d��O������`H���~^N�-u� �Ɠ��p	0�@p������>��X�by��`�c��� ���j��; ��\RQ)R�y�]�DH���~��Ɠ�M�D���׳-<%��D�½�����f+Ap|����rk���sbL�>06�N�\X�6^
��L��Nu��Ԅ�mu�V")�d-�DK�Zm��;�Q��n!�B�4��U~4�]/|7��[�^��XUm5���M�������Ӷ�:���ôw��i�g0�`n�m'�^�7Ts����+�Ұ�$� z��͢�4�?�ﰽ}��,b�o�R(�.�2�5�#��ד��j��fΏ��nC�W���6RZxs�\��Q�8�>�r;�\k�a���q|y6K�����
� ��хP��#�E-8S�,C9c鴴8:m��DR@�q+a&;�v�`>��|�����b� �Dᴝwj)�v9�㻱�#?s��g��^r��]���C�%caɑ3IO����4�G��W�~|����N�IEnADP��g��6�e�{ZF�lߒ&ҳ|�	��sj�V��"�&3~gK�&�~��i����X�:��͡������@�����$��)��������R�R���O�3�&ũ������eĉ�<����O�0B���?t���
2�V�{��_�T�F�� '��l󃂴���O�{��1Kw���=���q&<� ��+w6#aǸI���\��LL!*�x�<
V��ͼ���(�`IYl/�̄���o�[�����tY����������n�,g=��|ƤSY�"�^��$e�E��
k�:���B�3~��"�3@��X:��ot�WӘэ~�e'Os��B�~�H�����9�
�����-N��\Q�P�c��M��I�/S��茆�b�`�b��q'�s��}�Lu��z��yy���_x}bg%�}�u!6�4�}d%|mx���L~��K9 s�����GII�����m�"r^�g�{䠯��;���T��XZC�6�o@h$M�7 �����k�i����O��k�@�`L<��*x���
b�}h�� �^W0&�l a?#��/Q��G����1�Ҥ{��)I�׵��e�9�ϊj>�I ڲoܙ�#��Z
��:���#�p��\!���v(�_�\�/h�/�3+|xr��s����D��H�����!�
����ˏ��3l1=M���0^Mj��Q���֗'�}/�����K��
g0Π�\~�Ћ �w��%/��GO��-0
�7OV�p;�����k�6�׵8��[w΢�T'y��V�"�*<�����%�&1i����y�VN�%�(�F"�
��v�v�"<�c���!��<FJn�_��W��[��47���g��r�؍�e/�v�E/]�W����~\�9��CO�\4�,�O�-�� �l�z�̱DnS�'�U�;��j���9�A:S}8�U��24|�<���un^v쾺8��ا�0���͛K�*8����e�瞬�Y8z�=}¡�w��s�24�n,>�C��m�m<o�����r9�R���,���8O��{��c�|�0��4v/���ɥ�3�Ǡ�d�����N��܊�\t�A����Ȓ;wҸk�4Uw��Χc��]?c�����`�����Y��H��.�^Pn ��k���L�p�L�R
S���j�R覀u������Q�Ã�(�Vtx�,T�T���
�z6 }�BރqQ�]��1y������bbc��L^�`a����@��{9� ��:�U\��'����F��I�H��ϙ�S͔�����l�y��R��%�3*�m�������c6�'��8! ޻︬_��?���k|���,�����_�MV��=Û����ÂO�9��$\���U��_j�iw�xO(���Z`�<��h��{$2��B:m�;�Ps��ĸ��i>�|��V�� s=M���-�{�Wb���B�YA��`�PXZ�W
(؆W���
E�� �(ڀV
�j�vd�l�"�l�G�X�'�~Ȋ�J�8)���{ {b�����8��v?i��z��e��GV�3�z>�����h_:%�m�M7�BH$�R<�3 ��l��1��i�y�X�ƨ���;>�=/���1� �J���CⰟD*lf]���T1�0:aY.��2 L��HRiG���4�|�^֋�l8^��n'y���׊Vk� ��G�+7>F�����c�\JA�����@�gkYʚ2���,��h)k����yBVwp��ȩ�$��aL���_W�l�s;%Y�)F��
� ��,J���t/09 I�J��c	~����	�Dd���e�g�J\������M�`��^��"��$l j~=�J���~��]H�Mˀ�QT�j1�3ƻ��L/i��픑�����!�s	��k��#ߧ
~��ې?�q'�]�L��c�#c�N]�=,Q�����8����ŏ%@�1g�>_��j����{s��W��"͒�*�S=#*T���`=#%|黯g'^z�$�%-;��*&^`��1V�toѝx��{~ƞɹ�Ȫ� UPSw-Ӈ:�[7��$��Ȩ>ݦ�����j(�oۚ���\��Ḑ
�� ���-~�٫���@��������N32ƶ#����A@~�>��o��)�,0$�$\�e�a��$�Ӻ��G�{�P~*m�$��
���d/��c��<�.;:7|"��Ƹ������L�~��~ؚj��V��BN�P��?�����e�6�Q��9��M��r.�#*/*Ø�'/%,-�l�-5	�M"�E����~���r��.)����fN����2���}�-�|��8(�$��ѡB]�`�l/�G���?ޅK�k�m��-�ܧ���x7��]+Df:���m��If���@pJ��s�K�� MrxVU�L�WZ@�P������bW��.Ƌ�v��?8���V#�n�m�A��~��	�d��M-?����$���Q-q}��ɱC����2P}Ӿc5t�y���ɚ��]XŤ]H�)|�I��Q g��9n��	��ͭrϴ�:��U�����O��9���������N����v�ļU&��v�@¢J-��w��EzO�~
�I_@0�J���ڃ~��M�W�IIE�~��ȍa������a;�nN���Io��/��[F�°B*�җ���S���?l��u�}0����(l-�fޑQ��3�`����^XF���|o��?#pZ��j2���d8�[������;���a��%�fR��{�C&���Qp}54W������{�:'���C��[%���.���b���Ǧ�a3�_#e�)Z$�&?�a��9Ā1��T�ۍL���z-���N��|�&=�,YK�Ș�!�9p!�<��B'	����g�ͧ��?,W6?- �c-�~7���Cig���m�g�D�>�3����j���Ho�4S�H�/�YwZ6\]��j(�L	�.L&�dh��xg�BT��@:ϕĜg*��I3x�h�a��|89j�)�ٰ�M�ԣ��ԣ߇���QV�O]k��F��*�JW�I�E�}?��8�7t�a�8v���@hD'�D��r�먶�е���u>|�|��̙{�Yl�B&ʜ����X�\5	��%�U?�Y�j�ɳE��W�"&�P���j�t �zD��z~�F`k���AZc+v6q��Uq��3d�خ����s������y����v�b�_�۾�t{C�{�sbJoC4
�����Jg�ҽ�^{��C��Q3d_z�V��!���p_S���[ O������{~�+�:;�3,��./.�&�F�͘�`�Sg�8233��|?Oے��ǖSI�hA�����D��� je!�Liͤ�KP_a��"�
�R���p&�Qɲ6]Ki5?�QY�ZrGRV&���K�|Sv�:��-O6���)��%�I{M;��tx�ΖİȻŎ�f�JIT�o&Z�>�L/F�����uFq�2�����@&���M���-f��F���f���oW���%;5��U�3�,�]]�/K�#=ب1�#$��i���v ����=�d�@�u2����(��hA&:�d�%0z�. ]A��jF�{�jd�0��ey�tyg��3�5+��MO��G�b2��(�ջ���R�,(��1�.
�t��X��������H��iP���t��O:@�+���r^z�����c�_��v�"pC���m%}wְ�/J�b�A��:�4��_ǢRh;�:<�1D #�ҵ@�`Gg�+��z�H\�Fkg��T
�ɫ�/E��?��3�Ԏ���+Z��ԘŌ����R���9^W}���51"ҚA����z;b�b�)j�e�ڏ�/��:�#�'�4{+�q��W�z�K�Pcҩ���2.��r{;k:͹�Z�5���8Jj~p��;��B��� (Sz������QTS�cs�Ы��{��LD��Y ��	���i�	�`+9��`ԙV⣸���e5㞋4,r�"�B�8���O�r��˭}�'_��W��@;�`5�S��ڥmh|L�Zp���46\�H�{H��p�� 9�702��z` �HG6�AZ*L�/ơ�i�YK=�щ�y�lH@�p�K��$<��t��R(b�/z��+�w%����U��.T���ӧ�HjGt�FL��*7>���C�M��S��^�6g�j�<�/�_�y��7��V�����A��j��ۗ��T*�wX-?��]��vC�&2j=����G���:69	h��sǎ�#z[��W~��׏i�����]$Q����U�yIk�t�g���� H�SE\#�_����4�j�	�[V ����ݎ?�8�z[�w[/UX쌝��3��Ĩ梹��G!�	��T�(��{;�
�>D�VY��������|��q�M:
�{'1�,k5M*_�%|��ä�N�ч�w�֝�PͫJm�?:k�w��(]����߀DX%)g�;JeS�]���W��EB�lLM1$!�v�*䳲l�:���}m^���ՍX��i���.���1w�a	G�4�U���p�$�2*�~ƯP�7��=��qđ�=ĴGA�r�<Შu�����Jq�n���]�\�,|����	�&�eQU�+���_�k�ێ�l@ZĻ1����p�/b�[�@�7r)�; ! ��A�i�UM�,⺡! �c#܆dطC�*�r�FO����~_>��9�4�"oy�r��$��7k��颩|CV02�����;���x(i���%N�4��2c=pf�!U� �N4O��ׯJ�ʻ�mW�dA8�0Ai�t��W�*B�f����]]��l��歠e��HJ��)So1��9J�m8��E�B� ѓ�hჀ�ꅐp�h�v�a���c.�T��^P���
1̠�-_4�]�n�Zk��P����M���K�搆l0d9d�P�����G����y�,E*��	�G��m$�y�Eq���7���D[)6�U< �� �:Ώ��k��X���3�g�#����X�ҭ��G�E�	��ʽ3�`���Ez�M�t�X
����$�3�M����w��oN��o8��%�0���TS⣍8�����k0���x���R�(@-����SQ�׬]�_Cܲ��'tU5�{�<,BPFN7��$k�n��JC+�q��P�Y0�^���)���Ef$�Ti��D�xI�֦�$��� �dau�� NK��,Opj �xyl���鲑1O��ҋ�)�'���g��*5R �d�Q/�H���m��G{&� I�_6d�#9)Qys�j�m$��{����k-	�̂�p�?�vXKG�K��O:(�' ��e�'2�OjU.�D��Д�&��g��:]��ڔp٦�Yއ��]��%\'߾��nö��$���wJ��pt[G��"F�EJP�ߘr�]n�k���JM�����9��퀦�I�@�+BA!��Q���������[���R[7��\kf�u/x�Ko��`����R'����}��HHZ�dD�Z��R���7»J��/4dǏ�����9nK�����$��ߌu,�,8�5�. �jzq�[8��P�2�5J���ԁ(��xTQNp�Z��)�R
��!�m��l��<�)<�X���	
�Lw�x�K���"�fQ[5�BS6�V��2}�rvx�#v�2��Bd���U�����Q/�[�h���X�f/�1qzI]{ℑ�+-��[�XM���$7l��'f_�y�A���#D��3hD�YQI�8 ]x�s���j+tY���#��*:�U+k)��S;߃9Ŧ�kh+�	�tld믕�BG�	��Gf��q��|��A�+wi��!���=S�E����B�����E��i�S-K,
��f<�����F��V���S��cb��Ҥp�������&ϾZ��y��2�ٯ����Gx���������� f��G�nPu�Y�F���4Ҳo	���8rU�d5��2�֢x��"A�v7L2��œ`?P�s"81��Ҷ|6�/��5B3x�!r��Wf1����#*��<Wlꉂ���U<޶�H����F�}N�iA��Z!�g�ȓ]��7ک�9 !�I"���I۠�p"�HI �^�8?ܻ��,?3���uDڦ�vL�M�h���q|�D�]���SK��|[��"�:��+�ʔ���t�e�"���P�����aw.Y6-Φ�\^´������-���UyR��^�5����h��c�g!w��P��t���ب�6�(�CM4Ju=��iu^�����A���[QƯ.�&���k��������w(pay�a��Aլ�0?Ƭ�O����0ᩧ���g��>�G�م��9&��)���[��ۃ�=	\1-�<]������9�ܔL�_O�i��J��sޛ}��%_�'��Q5³��_�D��V!���bV�|�}��ߪ�Ep���i���&�ozWE�]E�f3ܚ:��\�Y�H8Kx��?���.hb^�,��ɡ�R�S���}tv��	D-��7��a�}X4����d^���^�y]pr���Go|�RQ�z��)#WjlR��R~�R�}'r}7tp�d������U��{,_C�CD�����?��P��?Zq��3��� �nN�AX���&h�PȸҢ���J|�p^�Z��7�=���|�g6>��I��>��we����I���`�J;C�.Z�)xnv��3d��q��ø*i�9HQ����ʟ��QfFR��齆dyW�,�2���P�ќ��=��fqXv����v�<9���U_~�S�=8���� ��̦��v��X���t:����LG#�34Q�!����5_�N�j\�i`')����
R.��2���&����?~!�_T^�f�]�����}�l�_�K��<�����a������tZ���?�F��j0.��t�R�gP�A��G`�҆��p�6���/rO;��O�ZX!YG�0�y�O�]�3S� qiآ�<1�j��4�wD�ʭ)N)��>=R"����7zS�O�Zd��\���ի����Q�m�,�/��X��� ��'A ���9O=<��i���}?ۂ��� ��7U��[�~A�Kn��%K���v���#]�Y�?�;�Nˍ���,u�A54!��Z��A-�����`3`�'�1��@�m���G�v�O��p�fQ���[���صW
f�6��=�)�_9��q�����Z')�lf�p�N��t�Q���4=�^ɪߩ��/��'
94�϶��1�M��/C�����RF�ħ���s�����HAΊQ���ڢ"u��m����qQ�z�r���`���OJ��ꔈ��Y4��T�YGm���E#!l��Z+�uS����e�>m;'�	��ܬ>�E�̎(^i��Զ��P�:Ct�Q�H�G�L�������5��������k�"�4+K%C�k�z�(�-��mp:�a�@���<�@,��ajm
��K�Ü�>t Y��]�qȊ��}x�E.�<0>��l��X6���|$.މ,�O x��DC�M����ʀ�AS�Í�ds���"���by-R��<�^C��JDӈ^6���[���D�x��whn�Dx`T�x�̑8W���W�4�<�\%Q<�H�Z;ed�l|�?)�T<�=�UF��4:\��m��Ԕ�$�	�Df5���=��u��Q/�I�����vX76�آ����7�q�ѹ��rEѷi�b��`Ao��.�x��5����-}�h�G��M�nf�-^���ڴ����x�8������1�Y�)��Ȋ��s]Fw���y�P�0֠�1~y	qǸ�uu+�*�ϩ�px|�u*QS�! :�lԅ�0���5���\�r"���WZ2غ�����7}U�Jb�\q��R�)щW�t��L)j��f��r��)�%���#}�/QB���MX$��I��v�~s�����{�R֬���˔NW/l��_޽��ǘ�Fn�5��Y�����_c�[�nY�[�Z�������	��Q4S����coB=/9�JX���SCw
�fu>�
v0�SHM�o�xqU�U�Gy�����y��`���Mb�x�߭ �_�o�V�dҤ̡e n�YoOT�3��ל&��3k�+�c$	��~]�f���=v����wŦ� 6�b{� (�����$W�V����Z����*(A�B�������ų$J9�M��9���:�����m `�M��;D@D�k�^��зu�:�ñ�x�G��7��Y�Ֆ4pU���)7�~��@����f&�H3n
)�Ku�*t��I�_k
�#�7�^���q݇�Y��׎��������=f�������jf��SpQ
v�[PF�(�Ka���I�XWxh��Yi����D�� �������g���@��E4o��0�tz�A�F;�V�Z��U�p��f�����aQv���P7y�`�M\K� L�p�J^�]h����Ȍ�b��CQLm]�*�2)�(�Vh���LQo��_���!�3���L��[�_�X��@��(�n�y�N���{����^�|�hP�.��f+�i"�������'��=�	 +H��͇&_5���kŗ%��%aV�B�~�kߦ�Cl9'���~f�!ж�2G�?�J��q�M_��h{�*�kW���O�L9+��z��V�lτ:��]���{�"�m,YA+��b����0��$Cq~��W�3�?d�_+�n�
ϯ��K�?�hq���C�l�D�>� ����Ҫ8���'��G��p�YӾm�����P��� ��w�Z6B�֒m�F�F�8�1u5��%����+.?T�?��<�X8|M�CW��>��k"�)Rʖn{�Z�G��h'�N����x�)&��8k���r�)dXuĎ���q�]>���>dy�E�,mP�f��żO�ꑭ��_�c��QK�&r� ��i?+�S0�����rY��[�eAj�g�8v��6�������@V�� su��p����B2�K�܂�i�)���%���փG��Cso�Hr�|m�ݱ]R��|�ۖ�M�Ս�}��-�c15�g���c�m�Eh�͟	-��/�d�8�zp*Q�@3�8�6F���Ͼ)R��K�4@��]1�5���F��㴵t�f��vr� 4Մ���4�.V��W�}�pǪ�z�	+q5�$�H"F%K�ro��$PN����E�+A�`mn(�ka˻�`�ـ޵��}�=�'��x89�:Z�l����[��\#%SQ�M�(6�����N!oi��'^r�
��$�i�<̗"���T'O�	!��Ї���REʘ�~Q�!	�,uZEt��t`�=�Y�7����v��C�2��l�F�_�A�s�fD�y�9�
�	�[���fژ#�}g������BH�-�QԖ�/쨊��E�{y�� �!�Aj�a%z���8��M�>J��	�x7/k�z40�`�LWp�N/Tl���Xؙcܰ����8���"`��E_:�R(�R���N4��S-���=����-.�#���6^"�|��}�Ax1��2y�D���#�B#���{�TItr�bԵ�=�ox����4*nފD�Z¨n�7�M�q 0rҮ��y��)��Fb#��8�)G����P�;��-Jz�F�F��=�\�X������E0���`4�G��u�#�hZ��G���Z2���>g�jv�4xY�!8�ۍ�;߰�
Uz6Yɋ�DZT��2���G�t��u�A	�k{�����>��|�PP�c��Վ{�.!KL+�r<y��tVgg}5{���d��(�Q�m5����;|S��
��A�jL
5��1����JA��H���4�! 0��e3|��0����7��:8���&�}g�:�e�x_]�gq� ٟ�Q��U'����!޲���� ˧?��c��ܳ��Y��d�h�
31���VQ4�����Q7�!&��'|ֻ�\��O����/���Ib��c)͹{��^N�SG���$���f�q6ԾE�S'������UcK�=���oK�ʴL��w�!�p�O��<��� �>i����f�	���A�����ħ��
��haؕ�-t`;�幟���Y�uE�kD �K�܏��~�H�qV��
"���%��j�*%s�>_�q�.���2S��B�C�S�앦��ud�+��α�h�����Μ�Ō�D�����.���M�/��(̙��xHwCH���5����Z	�NΏ�c�J?�YXLW�xߏ�
8C�g���T!��	��k_N�oF��P��+�p�9 �Dp�`ræEJ���I��ϙ��zlqLI56a*�B���k݋���@�����=73��1�|��fL\����([�����2�o�6u���f,�e^�F㶆�Fn�-��[jy�1�2L�$�i0�"h�ܯ��}�]R�N|zn%�]]� ��'��z�q0�5"�h��=���*��./��e�k �����"LP0��Yd�Lv��́*a��Is�b��q��o��;<�pg"EE�����\3�6�=0+�D!��~��iۈeؾ������c5	*�,h uq�_��L$5Z�xU�eA��"<��9x�Mf�8>#\]�@ƾMO���I��� ~�bȋ�T#��)�A��KQ`���~-���B���z+|9v5@AZ������9�'ݲ3��z��Z��P���`׃����S�Y��t@b@�Y:���Ok;���0���*IBG'�_���s���I�v��`�,��ſZ�_ ͈u�Y{+�6��Qi�g���u��WnC~���\)�3CuJ���R��[og*�	D�I}���`�?濪"N�*|�nIx���&S/�|�RW>m�wR��i�x3��e��������[���X�Ӓf��t1��h�����h}�6M��%mT�7�<���gXZ!�6���}�U�����ًo��-����}��/wNH���'6�t���D�^�ta���s��r�5��E<�}^�O~t����nPf��w^:^�N�m��ῳm`(kj��h�;S����3��k�y^U'1^Vg�P�X��O���u��/CoMS�Io�Ɨ�l@n!M�	���nG�o�I��gD8e�;�-�G[g2�C��t9�n!�g?���♢�w=�,G򸊣@��~q����χud��)�:��2R��F�b�AV7v�YF��x�V��ص�A#�cKK��D'_�R�g�G�M�p� ��?���w�d�6mΪM�g������Zv�43�"gkXk�÷���,����ZM}��-Z�w�,���fJ&%qk�K�!v��o  �����i��7t�[/��ބ�9�"����k����ږ���L�1�Iڔd2sT~Ш�Ӽ�}1im�{*%��0��f���>�wBY�=ǎ�[!�?ua$���LZ��PJ�"��W&��C]�W?�o6������Ǹ����r/)q	,�ns���a$� .�E'��0kO���̵�3H���g�cNo5ڕ�D��%"@�=�Vl\�.���{�7uV�.��gC��I����v搉�X���u�/�4S����z����f?n�۱Aw*�$6M�Y�T�/c��/h�]'����D�X'���N�a򚽐)�A3� ��1p�E�f��nض�����m�� Yh1h�-ʨa�{}��)no��TS{���0���Un�`��_ͥ���z��ѽ9%��m�J�Bm�1L���V��3̌I�7�Z��>��u�#����[A�X6	<���-�$��i	�^u��0R��CJ[gU�'6���i��aWW���
���%�@�'O��Z"lo�V<H�]6a�o]�1�7_�bD�u�-�C�_[��2O���%m���^>�Y�������h�ɐ��=�x���U����	��w�ؓ�6�E��
]{>,:�lߛ�����ʨ����OcN�}365.�3MD�[|��[�Ӏ1�ؿ(ns�#pl��#�)��@Hx��b.N��_uʒ���޳NX)Z���B�NWD��dX 0�z�d�W�|I�T�]\3�:<c7���O�	]k(Hb ��� ��8�S�7��SYY�!n�+>&�]�"�X���F�\mG��+�b�T�g��E�yn�5
Zӆ����ũݚ����S�1��8Y�#�?P6���/�Ag���8�<3��7���9rYM�s㻔�\7�d�Sm6��x�z?e?��7�S����	.�)����h�����5�Gkm��^��3�Ԅ�dB����XnH��������Ԣ96ϼ�?  4@��3����G�!�԰�Z��_r���᫷C�������d��s,Q��7�����a)͗RZ�E��l�L�����2b�ꓘ)1 �vf���(S80��o�0n7���ʗ��j-�4Gnv��نn�(��l�Y��A�ߟ ���o�2$s�� 5}�]=e��GC�{f���	n���a�G�������	~�?!i�P�BP�因�膴ez7���I@j^6Z>Q���[�vL�|�*{g��H`۔"�Ș�w�M!�ߍD��P{&Bp��œt t����̜�W���:J�-փUb�v�s����P�����C���G�����Q�����.�Y�:y�q:��u4�GEq�ɒd��������S`�0�0�ǳ	׃�`~�C�t�5�Y�J."�y� @��_ڂ�. Ox){4����<�@�2�WK{��~6�T�C�`��5��7s0VTz���c=�|������|]�&�}U�[�Ȋ�e�z.�y�7��wK�>[�ڵ-&���[��u'��Ο4Y4+������-'m��_:���r�ȍA�<j��>��-�_��=�����<N��K��v/�B�L��(�n�$xǲ�~	�5WW\!ɂc��{�L���/���/��Ħ�Zr�Fm��^�y�`Ԟ�u� ���V4�ēe��)�.[�,�ArF�nm�lY^=�D�q�T��h�/��L����.�2LaUi�%ٵ��H���܆�vL��1-�@9�{Nt�b��ɻ����lf�������-�D&��$���$?����?�x�𛍎�;4�^޿P�fu�k��91Ɛiιk��bеټ�^�:x=)�S�a�Nq��,�o�n`��_�L�\`����u>�֍���x�������b�J9 /�b���F��Y��Z�Ӌ[�	 �^�ލ��^�0c�����S-&T��ᄔ�/?�ms����>C$�MU��K`C6�Z��7�v�^����
�]�}���ی������d�Џ�*xţ�^j[ Tqy:w��_�~R�3@��	v0� �$���x�G���%�$A��x'��W��o�;!������B+��\����w�޽PB�����9�Jʂ�cۧl,F��Gw�⤡�u�%RɌv�r�A���S>B���N<�����!O��J�T*��+k��~�[�����
SU�ߞE *I���N��k!!H��B��N]m�Jp�`īd%h���W�cs�2)j2��� (G�Od����:x�#Nk#$���VU��)WW�;��P�s�z���
I<�$_�����<��d��܎6���X_~��D�۴\�=��F�c<T9���֔�/Ҝ�9����s'���|,��/���x���壨���iRV�3L��t����!���a�~£���GM 	/�t�:M�����p
@&���|����UG�0Kܑ|�-����Ob\�C�f�8*�o�
���%�W�G��e� ����u%b���ٸk��Ɉ�]r�ʽ�=�/.۳���-׎��:��wqw�PR��}�(���A���K<�:X�
�Y��<�,���[:׏����X��N�RV���:��3&�x����>hn���:�z���˲O���I+��Sl!�\)
lH��<�V>�S���u\�륽�q-��������I�u~t{�� �b�1~>�c� kՠ�)��
�}A	�>�Y������Ly����|�[��X,}�V�^��i4�]n(�d�׳�q��O!��ʼ�cD�Ql���8tP5�G�3�i�ޮ�;e��W�\�܂*/���L�U+o��
P��Q૖�?<4
�*Z��"3�-����P�����t]����]�_�{���Uy�t��;ں~�󊹄f4��O0C��k7m���؏	�Ca�U6��>.�p`�R>Gxz��i��vac��jk�,5� ��#�{�D��Ѹ}�m9�P��4�7�ģ)-G_h�P��D�H�Yi�r���Hx�ۘ�9�ˎ��IssϞ��Ҵ�N�����x�}�
�H�8����<c)'�	l�G���Ő�<���O��9,q&W�$��k���V5�+Jѳ�k+�e%�����8G�N��T��6�l���0>��9Չ��5Y�v!�VR۲�<�m�����^��QpNA�о�֐ׅ�os��QiSQ��~���]Qª���
]j���##瞏���cد�q'h���iV�Q��"��F�XΒU�F� �76���Æ���V�Y�+�]����c���/�26��ʾS�VS�'tI	a]WM�<�`�� �aFBs�Q���LL�ܽ�z<q?�IX��~Es Ռ�i���A��S)�Q�;e��:�ڶ���G��H O~�O�ƀ�����ó��Y��9qǋV!���v�
�heQ�۲8N���D�B�+
��� �!ȁ��g0ɜw��AֈZA#�D��u��o��N�C� ���w]<��Sc�:��;*Д��N�)����6v� 7A�uumFH�@����v��{�iڤ�6�qm�5��J�Ŭ�XX��~�@5j\�2vso��#轃��w��yiR�,fI6�~G��M���� =���v���x^���%z̐����(%�b�.��p+�#�GݗI�+声��h���S[8m���\��^x���s2 v�I�?�hLu�\M�]�c���@o�#>a��=,>�6�nPѪu;C�ۡ��j�7���!��<�;y���<�V��儈ai��O��� �|g��<o�m�ZR�����ЖYJ��r����{���;��k�.^���J(S�u8u,^��6)��bt3��e@9�
�a�>ri��WE�k�ܡ�.�C�tb�C�����\��9�2��N>"v�@�-#T+�[�����vqNs�5N%m��t$�6#	ɇ#�H���e�?u�J�F��x�7(B��#<
͝Q���ͳX}�1f�{�2<����555���F盟��;�!����J�Mi��T�v���V�����ǿ��$u��N�˚Q��%NQ���TG�`�}f�T����]i󆫊ah�Y��@��|�eq�-DG/gzK82�\f�9ێZ�w��ɿ�sW�LU����;A&s�,�+%��{ L���1���P|s{q�n	_���?�]g8�/���3����/`�alR����~�����KƋ /��3��:�V��al�Х�:�6j�c�ȏ��ox����T�+�c1�w�� CL����5G�0k0���$�����o2�=<v!0_���8&�D]
��YP)X��E{�&��x�1>�u�d��5]�N-��=n���im����H�����G���|ܑ-�Q��'�7������cjh;��Y�HNZ�7������3�|�>Ĵ�~���>bq�<��b� l_]l�h�S�Y�|�os�L��W��V�h*�f�/�1�=5�8n���F�\vW�)���F6��}�׮�:H]���kD�d|��
"wS�e�~�5&m�&����+��3BE}�!�� ܋Kp�9v!=0�e|[�1���E�J��@�k�_�pE�|!NT� ��?&�~��,`�ӯ��|�3��>4S�Z	8��������s˾��_w�U?}-�
T?�b'�`^ET|��%H�|K��lw�f%���Ӕ���R���ΐ���~)H��s$U���IfeA��2�Mk|�r�=�����vJ�ĺ)�c}K�#�ʀ	g��]�
Q0�c��}x+�t�e.G}4��pj4o��)+,`^�[�>�	k��)���Ȣ�7����ᷙF��FxQjҏwcd�{���aN�\�f��0c�D�%|8�Q�X�hB�[��=Z/��30W������!O��6~zU�_���j�2[jx���W� �L��q�q�p�&��dW�u�a��c�{��캒cH�Uc�`�V�Wh�p�pG@�,^��	����� ~�8����?H�(���Fh����?o�y��gti3�m���V��Nu��%�6����L��$������]|�@�8���1j<�D�[k�kS,Hl�[���!q�N	���.��pW:Є����샭�����ekN��q-�S3�rf͛d��81�X��Nx]��Hjӂ­��'ס�LV^�-o ;��$b(��(�I\��w�����;�z}�&�٠ہ��=��X�Q9I���x�*^Y��W�7�r��g�1�����'�8Ǐr�W$쓄���Q]�u�m�):2���%:�M�G�p�~�\Qr�T�Ę��@Ӽ�+�QoV벵��<�����D�8�|�K7��H�t\�#˲R���;�o@�X����za���bm6R��M�����nb��E`� ���@/($G�j��5*<�����x:��>��i�ub�1Tc��Yv_�`�E�8�?��ɞ��cܢ�q�^�w7��ZT��U���+en��b�Y���}���.y���۽��՘�^�qX4�ah�j�F�h��p#b�B�i����sA��}H&kH3:5��0�l�3��UV¥5��t.�1���~@���~�h��:ʽ�I�¯�|孙���.�{f��$��5�	�v?j��ǩV�;�FW(&x���
�bY��'���!򱲗����%�o�K'��j���ʝ�7��-S	�-]�*��6�;),n�!���ȑC.�� $����{�x!� �z�� O,,r��!���v����{>���繕u�T��yG�%
`=G��K(��.x\dSj�-j�%X��V�M�?X��~��XC*R��z
�}[|[c���g����yҁ�m��p��l!�L�qg�=f"k�wG)a�s%�WD"�ˏ�[U�m�!Dȩ}5��2�58D�������̸C9%�j(�2[�2���ٜ�Ң�5 j�T1ĳ������f���?����ѯ�-T�e8z.y�)[4�Q 3��_����R�a�gӐ�j�8�D�ɉ"�-0��f?��w��8ܗ���1XWlwߚ�+��2:K�k WW�n)�'�����P>���,ű� �������� �7�M��Y���Go����[�+@���̩�������}$�G�p�� H�X�T����6r	;d��pAJJq��^>�=g���
iš��1	�+�$V�ȳ%�<Db�&ή�>C�¨1���}��~В|�	��^2w`v"��b{�'7��?�|����؇*W�5@�wg�eq~1Q�a�\3����?�#qb����8j�{qG���� �Wei5.��X��R�!j�G�:}������ys4�J�M2u�a
*��w�]���f	�q�xa�
)U�4j��,��d�/�s���%����*��F?��a�nDj+h��緇"��:�֘��<�P�k"���|,��Q鮐]X�b˜�m�<G1�D�/e�"b{��﨤Kq�h����G�?��������a�\��S�Ӄw��rY��K��V{���6rj�.͒�(D$`��z�*$QH,�z4�p�b�������X�����<:<!�W�pb|U��[}�폋EqG
��m��3�H�$����G;��@<
�{à��U8�c���|l��^\Nb2��Z���b%@��h���[^&l7� �)��"TW�wv #�͑�
ɈS�~��T�Y9����Rz�ᦂ#��������/�1Nd��eX���h��M&����qi,���k0�&<0�Z �RYu�[�A%5�M�3��R���GH3����d���*I=)G�A�Ĵ8BOf���Nl8��4d��h_1;&Vғ��j�����6AP�b\�Qڬ���7 Q0>r���Cp�_�LEX]Ǟe	�V�y�n���|��T���
��z�5�H�Ƕ��uVsF�G���mv�װP^z�%����GQ�@=�a3}6�H�ly��!<���,(����R����k�%Z��N0���!e�&��6�v)x�&Q���d�n�< �v���]�e�61L=﫳wS�_�����DF�1��z�s�+������{�@ʫy����V���Wev��^���I��Xg3u�`W9�Y�vRy{�ݹH,Z��M�4�������4�߰�|(X������h�|ծ�`�5lV/�R�(�J��P��{���έ�����cޏ�.�F��z�oY3jO����}_�|�t�R*4u����(��"G��8��A��g�[i�à�R�C ��Đr[tJ n)�����<̮�*ߵ��ڋ̶�;�j��
��}��U�AkzS��1��a����iY�v��!HCR����L��
b*u�{���Wi���DAֳ������
9u�f���Qd�W���߱ddneZ�C��U��p�,?����	���X]׌�ϪW��lL� �,E��H8�X���lW��'���*�Ç�#3��~��f:�=3[t�/q���v� CQ�~�/e�O�u�l����Ձ{OQ{-��#�͘��SR�IV�1WN�߀n��rj1�$Ԯ��F��M	r݂N�u����'ءɋ���ߚ��'�	�	��.Kx iwo�����h]:��(�S%�I��rxD�����T���d�o�'�:��ۨv�f��F"t���c(*�r���s(
+mߐ�p�AO�ޒUDV�����"��t�L��Y��$]��������k)S����O'[(�jQQ�x҆�
~Fb���XK��L)V�C�?��M+�����ɸi-�&���O[q���9
�I�z��lE�0J�@u������:�����L�g�r�KnwN[�_o��HW�΂��haJ!���Mn���4lB���΁���D~�����+�T��0��($t�c�2E^�Jf
bY�H�H6�o�K��ʹ%I�G�K/�?8!\|`��\�BRA���|1gq�̲:��Nk/����cʦ輑3P�ec�Ф�v@�{C��=�y��A�����;(2��nE�[y��f����eBB�ȶz�tr�+�V ���� �;�3��,2��-���aF�e9y�b��sL�έ����F&�7`ti����.P��'��ab:���L�gɏ�]|ް-��)jB�i�	R�gT������ݘ�("��*�%�L��?/�76�xj��O�<̍�HK75=�����#|�uR�{�N��ro�S���^m٢�4Fꄏ�j �]a��qZUU.����`��1\�<h���b��A� q���{�@{�s��x�L�򞚘��q������&B%���cN	$�|�6q�$_xlin`�>�ǟ�.��{�;H� _�+/�����|�M��qÝ���3�������ȉ!9͐?��cm�̒�..��O�-��q+3�5Z�N�V�d�U;�q�f܋�g{?�g��i�2k��[�wF�yc�����{Ϥ\��;��d�ҩ���V��_���(lIF��r)ΰ��4d�!h��L eB5���F��Һ��G�T^�yKB�M�X^0���Ʊ�E<�"����fԇD�,]���x���P��~��`2�E�v��Ԋ�a0�V��^h���)��앍d(m*�+�A3���Ӹ�˚�xnwK��n�N'����x$����g�υ	p��u A��M-2�'����K+� <*wj j���*��Va"xQd�N��&�h�,�"�`w��h`�[)�u:��;! &U˕�3�b�B`�
xy�e5�U C��<���Q^����p�<I1Pr�s���c���U>�ŧ����g�~�\�2�?V�M@�{���!�ɽ��9xnYD=L���l��"���E�'��-��@~PM��;�q�k�������y=Fu�BߠRn�!�	Kp5�������
�c�^2v��M�{� ^6~�͊ؗ�^�w�.������e��+���:Z=zwͱ)��v�/诒	-�@Oٸ��U�<��m�����TM��,#��Mк�:��+L&���v�|�H9)��#�V[ùw�L[�+/�K�)9{�[;�˄�v��.���nq\ 8p���;'��x��hn�v,���h��R�M��ֆ��e#Þ�;)Y����F�u(;x+9ƭ���Q�&�q�үAk��	��ʦ�s��J"0�D5��W�$&7��I6�5u&�N]����蝯Ge��`�m��-��0{eb�"8%\<q��<�d��'���S�򨗤�*���&SzfrU.�O�8w����p�����!,}Z��K�1�9WP�QC'$�����7 ���j�R��D�NK�k��ʤ�,�S�y<�6c��5t�����-V��s	I����a�v�QF$�gΖ�4=3GG>��!�ѥ�i�"KUH��#�񇸟�
�q��[2,��-2�9���9 ��:��sRAU ����*�}2Q3�|N|,Uxv�1[�?4�y*鞉���""-r�����(x�>-u��Ȃ��_n;�	�����#>t#F@	N
3`�ǳ/�a���ga`�ղ�`ᗋgj=�)-�5����7���4�Q��b�LF��w��b��\eG��%�Y����gi{�]Iv��h��$�BSAL���W�1�ƴ��A_��@M}�L��?-C��b�F��&Ӟ�ig_Bg�q���p�y���&wD�zH|<��o���@0S�DXYz�r<nL�ΐ�X��(��,1���U��[��Nt8�uZF���k4���O�sJO\����@X�y�j��`(��=(��_]G���gP��<>F�.��[0��ϑ�%�#5k����ީ��EG���Hk.����0�-Y���PD��-t��|�6�g;H^X��}o�n��S(����з|�S_"[K(������{3���2��-8��AGpC�_���bx�?��-H�6Fe����#<���el�!�l�^5#<=@NR���~.)+�/���8�
'��X{�V��}\�S���۰{Q����.3;���J�8`?,1G��)�y�x�0�h��r�:,	�����3x���0���d|r���s�[ �����ҳQ�4H_B,l�\��R��sQ��9�-kDf�ܩ��r��ɗJX"��b5�V�p�yb.&·F
���if{.�=���!�.�PN�&�n�(%"^�qQ"�/H����\�(���Y�=.�����g�+����x������X�YM��~b�2��3��3�����ͤ�GL"S{y�;�f-<O� ��RӺ{�%�?$��/M��q�1�9�m���=�`秨����L���A��(F�`̶��QX�r_� �"`�#�t s
5��f�t4��z�E;�Z\p����B��q���3e��s��������#ٗi�����t��M�hݸiQ�0�ȮȖ>�	��A�AϮ�ѓH�O�� 8[�`�k�ھ^&�#
B�lt�x�Ecrf}P�'�x#�DP����ݲ�h.~�R,��0l�3��م3�.���+M�ʋ��r/&l���j_����tv%�Q�8s ��#�qm��y�hN�	�#G.���odR���'�A�'&���b��6
��&ˮSu&�%y��\�Z'a��1ܤ�����KVgf�����k�0�1ڏ��y�3��=l��b��9%9e(" ���E:\
;l�Fb%�<��i��h��s��ԟ}'	��?�)�"��9/:�?\������������1m����P>ӥ��ph�F7��'w�.L���5�.{��qk���6�g�;�cKQ|r����:yM���v-�u�<�0���/ω�#F8�瘾ʿ]X/�X����<b��K#�!#"��8��䯗}�0�אa�Ǐ��\�/�ZS��#�y�ӗm��k�"�Ҍ.�<��#�*=Nnܵ�v��[��Qm0�!���n�~	��
JS��+��_�4Y�t�'3���#��$Zؤ��ҳwf:�l~��&��1",ް؁y�Z�.�L:$�t+
�mK	!l���v(����j�4�AL��v`�2�a�;��PU��K�格,h�L<�C=���d��;<�-Y�Y�fR��x��a]�����@���e���C����q��|S��BZ��>���Z\MGV�h����&��Z����
��
<~��M���1a����6��M�n���I|)\�rԄ��ɼ*\�%J�O�u�W�}J~Lk�S	.}��_R�����h�o�ȥp직F�0WȂ��#*�U���_��w['����tq��٣�S�tz`�`���L���=�z����!�-Ks�V���9���te�` �}�m�#��Si���3!�VU����ǉ��n�E;�&�vP�� �7�q	�_�Đ	҅��hy����,������f����UA�����z�b[O�E�0sB��Vn�`a���;����x�;x�|�/|F�.қ�v�8�7�����3��ZY���|�G%m|��S�Ix���P1l�ArT���o�6���2z������6�-{Y��M�ou�}�ඒ��bmc��<i��tR�d�)W0_.�TS^�,����uk1xyX��i��3:
������?�v?��zFNB#޴РU�ǧU\Z��"X,��iL�� ��څ%߈ �����.<���N��23��h�?�Y�\���L��OV6P4�h3Z�U]L8���fJ����s)�z>>'���Uuc�����g������)� FH4�2���1x����;�]6�(�>Eˋj�TW���*�qa5��Wn
�Z��q��������Bm#�6���kA�Q�E�S}��B�L�gZ�J0�.VѮL,Z�;υ^�T���w�H% �4/����}����Ʋ�Ms0z�C�T��j��rm���w��ي?���m�<1 ~7��Te�h����l8�b�gk���}x��)����X�S����Ѳ�^X�f8UOF�D��^0�ةZ��!��Uy�q �=����݄G�Bq(���������%�y$��ǀU�����Ř��#�K6ء�6��>������7p�,�)Պ{����"h$x��_�*A߹��>����X��Ok,��������=k��:Tڗ3#Nގ���3������Nn�/��oY'�w�7�2!:R.,�Z��!5C��X����f������ƌk[{�]�C?ȉ�s�v� ����<~�����Tfs��g�����9In1}�ˁ���{a}�(]�N�������N�"�EG�]��f�%�4��L@�lԳGM��'T���n<��Ƚ"�LVL;_Bx_��)$���%s��v�?�8s�����Dd>~�<�g�	�s�¸�b��c�N��~y��9-��*յ��'����������*(����RW�m�~mg��/|v?E�f�k�HL��p���C�ǘBM�*�����䗺VՃ1$"K_��XV�]J��6�f��Z Q�<�[WW::%���QÀ+��+Y0	�3R��Vt�Jd��3��?� �ֶ�����Q�RH�o�Mg���Ȗ��0�hНX�Pk>�X���+��v�팁s 2��.y���S�	�F�i�D�<�2U� ڙ؄��;�\��؅�Qq�@������*��'� >��������d���`&�u�,��u�5*�@����H��<�;�|읾W��w���d�J�M��q�͡��(��8�9���͜��&�Ћ��䣮Ѿ#'�z+�x(��!��;�r�z�4�N0�.0W�7�R�Lj��L����>���!�p]J��i�!`�5(q�{v}�����@�sۉ�bf���\/<xcS���a�3�<�j�[�3�!��T�W�w�Eq+�ql��d�������6�o|j����]�|���D���(u�	/)5x��� O+���O�,���o�#�{��,��<�$�4����������@�I^h)��d�u/<�=ˆ2Q�X�=���H*a��W}�c!�*lWqN�B��!E<q���W鉪�a��jx�$R�j��3�������31�z�D���I�F0c����6H�>�> �U?ސeخ,���Ҙ|K��wX-������v��ߺ�n��'Pt�д�a�>��-�ôVp5��-�4Ï��v��+�d�]Ң�
�Hh>4����J?d&����'0�܃�_�qe�����fSy�_+�u;:\*���P�������YF�*]���f�:���sZ�c�ҽ&�r� ��v:�/�}^�{+��!�]Ѥ�4׷��%�>ML$ꗉ�� �V5�p6(����	-Ņ�ENZ��I��	!8n�$4�9���e�&T�27-"*�UxŶl�yY���!���-�Џă�QO�r<�YetMc[����(���$�����r��E�<�p5�P�	�x�!��X�~S*��ʽ�����߳��b��u?��)���^���O�s��b��@�ғ�����DVn��2SI1G7 O�I��^���S�l	�̯�
��dZ+o�1RӶ+C}��v����'~AJ�h�W4�ČΚʣE��DN�����ީ�6n�Zߤ��}ν��*s���WQ"�D�]H�?)�dTy���2(2�$,�wѲ���Ϻ5 R�(j��V�e���W��ؖǳ.���|�����pྒྷ�� �h��9�)�y��� �����N@��m-_
��{�u�b�ܭySH�;ᄒ�e�Y��:z{#?4fr�v<����@/
�ٟ7T�{������Y����d�%�Y����Ҧ�1A���_�g�sQ�j̐!g���I�S>����F8[gSi���������~�&�#����?��L����<s�!`�u�N���?��S��]{,';J��:H��[mmu��R��ј�/�V���Z�2���u.-Ҹʢ|�|���2��B����]�����=���eK"����n>�a䃎���ų�}3Y�!�Jkq~<M~5�J���5���]y��xXU�V��%�2?��>Nz��U�U:0o�y�q�L��z*f��'~��"��𘪠��?@L<X��a�vud@`�C<�	�K�F��S���U1��PD��=����4�&V�C!��r�W/A0���	T��E(C4-�K�
z�1Zn�����?�6,GNeKwg�̲_�ӿ�/�����!E�����0�?�G��5�`�H��m�K���}q�1�Č����&JRzs�5����d�OqԂ���{>rX��u�36��R�<�_�5�/����A���1V����oX�/2�,��������G��U�R,��,e .�)��a
��99]B�C�4$"��5Ω�P���{��xs��h���<e��Q�2��<%H� ����M��̗�U��@��p��k�����e���K����.a�'�m�Z �h��!����}�����O�s8���U�in�E; �^�?�ss.7ß����s~�D�KM<p1��n�:ɿ��&�}�S7�%�$�=x���^0��!��=Q�:q�������:���w:��kB���W+maS8k�F���swsCǁ��=X6ɬ �Nh`1�B�ĵ������H�dE���5w��0�u�\&�z���:q��ۃ�P�!6)[:�m?L�|��c���=�Zr�q�"7��֐,g���[�_0�����OSc�:[�y��%�lR��	�f��z�T����;� �@0�/����!�
q��&�g�0�Y�E��ŧ8{q�n,�,��;���9�M��|�)kE��A�j��R�CUB���� �w���Zp�O3�:�8͚��0ܥ�:��I������KUj*�T\�C�86(D�b��\��6GV������w����N�zh�9>��fK�*�* Q��*C:s�L�V+kwS]�ٯ�2�la�3��m�6�E/�X�=펂LKGDb|��t
��f�M�J�#i_��f�����r��H$�O{\YDE#$Y�Lh��"���v�86FJP���x*_�]���"b��mO�M��/m��\F�w��'EĆ�bV3�b���tp�/u��or�~|
��ڐ��?`>�\mI�r��y��4�9��e�=��$�1m3E2���II��z��??�my�Ewlq3ArT��	
�U`WI�lJ�v��k9�:8e�V�#N�*]�iT"">������yI;�b� B�����bԶ�1z"&�By�m!Eg�'��� ķ���x�@P�2�%�CL+�BN(�Ց: r��#�t� ��Yl����ōt#��;�f����gd�3sF�Uq�)�?�t,8ؒa}���kt5�s(���ħbf�0�&"�EyK\l��Ws�u\�l�
n�YZ����� SL��d��0N�˪���2e)љ
�T�*O^�Ԓ����2nt�Fh��e�.�i� {[���y��r ,-�C����rh}#{�'�e/���TJ�2�qC�w����)�>�[~K��HS�|V�Nw�<�a\J^tK��{��wߺI�X����Zҗ��K�!�� �d �Ø>xgg��g��?ӭx�̀�.�~r�]��B���<i�!�+�j��COǖJ��_�I�n�����^]Q`�dg�lcy}{o�3�6i	���\<u�%"��A@�xgqcǢQ����ݜ��� ����!�a	��nY�J]�A/�yxZ�����w�&m�u��W����Zs�J�(�0x����{܉��cR����v���.�Md c�)P8����^jH����E���ݫ�VV{��i�P���o��шuR3��۳���Q�%�5��x�>~�m�;9�����Gp�	���Y�mL�|�N�X.����Z��,���`9_�n=����� �����E�qڲ��ƙ�7�"�3T�$s`y�w�j�Ͳ$1>���q����F���AiS쟗�y�6�uQ[ou�x��ȅх��mZ�J{8\K��dT��IU�\W�̍��9��1'ſ�����5�[\.h���ET̏�,7��2��$�����XY�(�$�mA������r�86�O}^GM�[�%eEe̻C§�a~{8�wדa��$�gfy�c��:%�����ֈ�W�y�3�80?h��YIh۲��I�%'l8���p���)H�4a��9H_����8�n������G��/�)�N�u��n�4I��e�C�8|�6�x�t�� `��}�vtt[<+�@���9	�뷈�MT��d�w�0S�܄S�d��]��zƆ	z�`�$0a=�Ш}%on����ƼR;��]zڗ��Y��R�S��F�fy�Ę�vս�n���n q�q�S-�P;�$��ݞ᩽�F�#�fO�	6�ٳ��m
4�ޒ=�ъ7�-1v�Q���Qu?>��F�W�Ðp\e'XԷ����n��0�K̪�A�6�q�o����x�O��FJ
�#��`�}����:��-;����5q�uh.���i&%� mT6 �W�i�!:d�������&�Tܔ�|	x8�3�옠�t|�a����W=:���ٱ=��*.cl�\`��~�ڜ���]��0N$�Z!��+�4��N2 �$�E��ܿy �����QvHl���2��띴�y��a��S���{�G��Yn�C�&$D��S�������u�(���R�E���95��b��嗱@�1�Yܩ�����6X�+��J��F�gn�a?̔w���_P5��Y	�ԳY�R3�Sh�F�N�����c��R{�5ܾ'Z{'�T��|��w$
mP�����4�;{*�9��׬j�Y���*sqn`�V�!0�k�Q�a:� t�?�zl@혝|#������_ry��8�����K+S�\��ux,�U)d�>�rD��#<�]����t1����xKOX�(T>�`�ʼ.�]��j(���_Ů7{�\B��_����*�x��}�ӿi��ͣ�u�;5�lթ���-�,ז�s��{����������{6�3�Y�~�]�z�JDf!e)�j+�]�<fq7Ȓ�m�r�Q�e g�@0��}�:��c��lU�`��B�VM��zLy^+;@�ׇ����o�����B�^66l��˿���vX���S�^�uM��������X铕 ��/�N7���짳��7�m��w���b�_Tw�=zR�V�� k=)v��#Ո0w�Y\��9��>2"�UJ(��O
��u���'��h���7�΃��l�7�������͋���a`H~~�<�����˽��r�ꌘ|�fF:���������b<H=���h�(Y\��4�V�['Ww9�v-]�t�ل\�2��6M(~�_q�7�m��-9�e��$[�>��~�+���]�̢nRgb\��"Qm��rs��)�5�X^���=c[���P�t��
��m��dЈO����Dw�3z������q���9��7�6��cjʐJ@�� �`�Y&�8Xξ�>ls�y-��Gi���%W�gT-��G���r������N��󉈭F��� VbD3R{�[k~P�r�X�b&��}`q|�}5a3
�6�}w@�}�@>� Y���Ice0��%��$M{�����8��@��4"[�ذE�d�$�u�w�����k�����(�����B�]���h�7�����w�{e�rM�|�b[���b\&@bd4�}}�Y��/�>9�Qn�IL�"߇�]�zW�D%���ɾ�@j5k��Ӭ�G\��M,zl	Vj�r
��j1�$��lWcϘ'Z�8��di�D#މ_���� ����>�+���߉����k�G�t����thU���@���ڼ"
N���~D}�4�c���sͰ[�Q�s|�~D���u����=�<U
��,�+�K�j�Y�-ac��,z�7BG��Wc7�9�F��Yf�����,�(h��5�J���s��B�#Mu�r���w����=o#��~0�5��Q2$;u{ҍ~y=��=Ƙs� HXBv�O�Թ��DQ%?8���t5�c?&��9���ZRy�x�2B��ǘ�K��1�B�Yw$	�c=��u�K)�-f=`�kw���,9!�*W��!��B�{]&,g�"��X���i��yZ�n�X*'�p8O�!��������,,*�E~OEj��f�@�O�a,
��Sf����y)j�A�!�V�&�S�g;��9���ո�:��c���Pg��/��	dbl!�P�T%޸�����i�V��}0l/�dw(��H�n�ɵ*T�.(�Ь_�2m�,�g>i���޵�{��`�ʄ�ɩx��yB�ǜ�P���ړ��Uk��6�UP������T{�TYUD�(���l>���}iH���H��Ys��!�}���1}��)�J���R`��3)��C2Oc�x�ѭ�/�p��縏���E�(1^_K8�ZFS���>Q4VV�(�8��mx�m�
~:9v����!���M�ca��{��_��d�rV)WX�YIKH�W U����2����>��5e�R������q������3�����`�9�P�GJ!yI�9i��MV7�Rcj��S�̕i���a#:ġ}������`�J#�GT���ܒ�΅.����J�񁉠��n��sZ'?r����������~�n����=��Ui�ɑSVT	T�~��/!3� Mh
���!U�%_3����t0#��C5f6��Pp�@��dU���a_$��H۲@����N&�y!O���k�Y3��k4$��w��za�(�6����4:�~+Ԓ�>�\�A-���%D�>�[0_�F��lG%K�s�<�l��bk����xT����)y]���0�d�ۿ���
q���	�i��;\7ƅcN���u�
tEa/��w^u�Ȼ���6d�=��� 6���c
�u�m�����IyFmU�&�Ot��MI�-}~n��*6"�%M����8ǥ��x  ��u=��"u@H�zV�)/�ο�۽����L����B�����vFY����؃NOMk�$����N�ft|�٠Pǡ@�$#��zp�����di��y�MhK�������9�����@��L������T7��z����mZ�=�旞�X�6?�+X��?`��|��i1�E/�dk])St|17&�G*+J���WJa��H��8p>�]��P/L���FWQ��u<�+�(���`;��4W��|?��6�bi$��A��5zjCց��3GL�w}x e��@�%�P�h�;��b�]h�&w�c��fz6 @}l���4yl,se�5K�N�o�Q����}hi'�D�d|�5Z��џ=�������A$āZ�Ǧ�vҗ���c��`�c�ۮ��X�8���;hh��Iu�jd��� ���G�~
�sg�/���qqJ&��t��f%[��_Ur�K9�F�V63�>SJq��r�Ã�@j�VxmuT��b�AU<T�B�Vڮ���p)XC��<��A]��А�s��#� m2�hm�f��/�m�^ɹ]�Wü����3{x��H�ˏ;�:����K庌�1�u� z�����O��C�vR����g�{���"�=�����K�A��g�ߟ�&�4�J��.�ƹF>3hոFv�3 ��^$�|�ݼ�y���� 7pu 1��h�F��OB"��ȣ�O:��-;��!����%���P%vk�	�7K����i���K�ޠF��ƴ^��|px�	g�/�Y�$��݄�̈́b!�C�[O�D#�J0��ef2`��̼Tu�T�,�C��#��W�]<^E���n(�
>F|��߾�Yr&�ȖI�m
����ǝ����7�jR~���pv?���t5�>���akR���ZKY��!�J�'�u�A�;�P������S���t0���ܘ&���%���*���q/L��Qi���,�Qg�߽�SYR�yuǳ��a��w��&��G�������!9^s$��kv��q�)�(�ft�RP�~-xۉ�=y������;�
P�|��O�#A�'�5&"29ګ�z��ň��rO*)�+e��� ���3o�&�E,}����Fʷ�m�P�e�v}�ɏ5��]��6]uhq�Rܡ�+�������D/t�1=M�K�0����e�Ϛ�<uק_.v�����8���K��?���)�86���� �X��xU3t�r�gJ(�O�*"l�*!�K�x�
�f(�l����j�D#��@%���[�zݧB�����6�V�ǍXK�0 
�ؔ�ƝxCF��h$���J@,����m�*�)v��"���Ga�>?��AY젩:AaP���`�����_����JŃhd���������6�>�jD��dl�;D#��V昿��"���/�6 ���$���Io�/���|�>fU�	�/fOɚ>K�+��}���������R��2����'B�OpeT�'����XN��9_29����;�� �ˁ8Yɔ���2L��sVh�^(�V����R"ע�X�,�������Jk'�(��3d��>5(x3S���Hk�\�|���W)�hd�`�V�����ԟ-0����@*�,Ѯ)��z2Fe���S��&��������6��
=�>����α��}�)�',Y��>���z��F��ڼ/������]��R=����(N.$m�+����r�[e�S�J`xǂ��[���������D�n��o_��ɡ��a��(���7�;�Wb��Ȓ���8��]X�k���5#V�L�S��̏/��M����y��waF�谍U8���i��'�{ڽ:F=wW�u��&J�.I�1�.�C��bb��t΂��,@�U-7?��B�t��B9]�=�u.*"�K|[k����f�p�"��l�h���}�Q15�P7�����N�T'"�P�;�9�9�/� w^�L׸� ���v�~��R���&{�n~�#��E�&|!°�p`�n�����P�c!@|�C��x�'�ƀE��v{ʩ�{!���|� j���B�jy�4d��n$j�L�&��ϝSDv˷�-�d�h����(/Y;%�MW�#���~���^M��}�}�0ޘκ�<����q�%ve�c�Y��R�r�\��.t~KJ�����u�t(f���}O�xR6O�zB���������Aw�U�WA�0JKF[���I��ob��鞯l1��:1�'�$n ���F�"VY#K�I�~l�>�{�����������l)*x42����]��d�ΝǙ�ѽx�փ�j��h��َ��6����k�4�aIt9J�`�z�/<b�К���#�}>�$�SQ�5�c���]�9��3J��[�)�9�����U�i2�R���=� m.f�Iv�:Yꨠh�&Tq�.k��"�{����ő��y�V:A�S�
�=о��E9D[Uw)����7����.��DTJW��oX3�O`<���8�7M/ f���-)�q[]�t9h�AC�����J*i!<����zs��@x�[^�4�Vo��絵�׻��-�9�A��z��b�@S5��9�Y�`� ��G�Hw��gh>���Z��ALo�������J&-L�	3�u�N��]��D?�:�,�D�%R��@�[�bc�&-�l$k�E��U�j��1�-NQ������d��s�"ג������HoS�q�A8&���.	���G��z��m?'��둺���:��p���V�$�Ƴ:�H�"<�\)Sc���c��]�D�~�+��ۀn�it����(�쌽
o�Ƥ�u ����y]����@P8��W,����<��f̖��6�3sjx&�~_���R"����?z��W��̛��T�\ �&(�ߔ�m;H�vaJ�	˴'e����̢~̰$��tY���qິ��g"֢��0��D������+?����L.sd�k�]�
�c�$�ʑ�ǭ��۝�/��߮���j�r��~��؅�0�����B�|�H�\*�{���2��[��0j?ꭆ�3��,;��D�#kJ�(|��e8hR���o�ň�_ � �d�����R��(�}�ˣ�
�VU]n�Eأ�8+͎���x�'G���$:�XϯK'4.N��݀&kc����v�Y��[�KU<�z<D�\c��
L�	�r��TcY���*m2{��K=.�A�"��ݺց�����Ű�xF�����r�K�0���#����ڌ��&npy��n\C��1R}�o���3��|�����滤q�\���q���������s�ڋO��V߄�{
��!o�mK"���8@�-��W��k0�	K�շݛ�}��k=Ŀ��n=']�e���Td/&|�T���f�&U��x�6�ab^�/��E[�v�)}i�{�����]�x���ӝ�v`����8�>��8=�,����<
/�+�Y��:�o���dz�2�90	A*��L̉8�0|�������hb"��M26��dK�yQ<��`� ���`C!5��V1A��8�ťP�S�4�/^?zϵ��F�[�0��~*��i��C��7��KC�:¶� �A���{LBĞ�����y.>Bn~��7߸�!2ǉD��q[��7�F�jd`�]�e|����+��p�����aTm8�ȩ�=�R�<(��g��Ch ����>*;[�����Z�\�	���y655Ϊ$^@�O��t3A#&�i�;�2�3NJ/yE����+�+s�b�3C���N7ڬ*��c���_��Ǒa�bŧɞW�=��luB�q@S��>�n/[_�\-���όF`�8^1g�}A�O����@O��qX�kd���0�!���v`�Oo�B��vϴJ��U֙�7H_���cܪx��.�dJ;��ku���H�r�F|z��'ud���+�����|��|��"�@��x�~���؜�(e��M�'$[�d���7�)��,�77j:�1"��y���f���ed�K�����C�4Aӗ=�Ơ��9��� ���"��)�o9�s��y��@�dσ�h�b�	 �E$��rl��oē���ŷ��X4F������)�@��p	 (��<bz�}崯pI$�a$Q���-e���O#K��~�C��v�;�D� rHA0�G�z�~.�)�_���~�&i��p�}�i[��{��{�'-��K��pR�}&ν&>P�FU�\1��ԏ��?uj�I�#�H���[i����ʞ��I|���,�
!k�=¤�9ög�h�w�y �O���hlan������'w#<�a!�T�𻠆,��74Q��ז�G��a���!_/�Y�Ұ�Tw�g��0��J�i�^���t�&��R��{��},���s����"i�x�[x����ބ���Fv�U<8���#q���"���6	06;��9�[�%�,�^��d&�|P�}FQ(�i��J#,$�d�z9������5��L�Kv1E8��v_hT����!a=j��ǣ���n�����.���c��)�$x�R'���L�j�*V��.-���.�T�"��	����Rr���%�Kc$���Q����G�Q���VT�R�a�d}'R��]��i;�&���6t?����JT����H;,�����j�?�W0�s�ϓ��Q^c=<�(�\A����N�m2�3�s�Xg/6
&w�j��/����}��k�����B�9����j�f������&���Z��w_��4�9o��_br���}'C��R{�vߜ�Sk�Z7R~'O��P+f ��_~#HS�Mc�z29wI\��D��&M�S�4m0���_/���R�g�zک�R�С[���x�1i�H���Q�G~fOUU��3�V�D_�^�'��3.��Ϡ�ŁD��ך���KH�$��$���L��#�)b*L��e����J�F-U&xK�%*|��er`+q@'Cn�&nf;,;�-�TEj����������,}��8C*J�r4km̂U� E�s�S��YP��ǔ��Ã���~�v=�߳}�cm�X^�f">��y�FHr=T`�h�/���a��3h���(�jn���������PthD�
��>.@��O
��^�XOJ�����b����<&�F��7|2�k���. �f���u3f����&,��Av����)�7TȘ�\�ϐ�"q���d�J�*���x(s�J��tU�5Mr=E[���3;0��	p�a��,+rց�QA�o!�ƫ?�}yp�$������ ��SD�֜��MGs��Z�'u�%��m��Aþ�ª���Kku�� 
��r�~��Ĥ����A<O�*61Z�`a�J <m؎�"0J�.�BB���d�o|I��ڡm�y�)��gs�^|SI�V��a��1}�KzvcP��_}����h9����Q�N��Mf��[�'�}h�E���{���o`b���Q뇆�3Jap̉5oH�������֐7�o�����<��}=����`a{�Բ힟o�x����ӗ��!Z��[o����pD����{Ú�9͝,����L�\
?|�ds��C(?8�7h�D��<��Ä�������'ۖ����~F
`V��>:�2e�m��}����V��p���f�U�sm�d곭��ׅ��"�\
&��N�0��g��Q��qڿ��D�]����]b�T��B�5t�Y.v��]pzŋ��m;3�$����VR�S��KK��x���韢�8/��EME׍��W��P>��? �0rV��w]�%k��r���:#/8��ݍy�1��c �@Z�7s���0j�7�P"�yx�����Z{}�,�[�]\u� ��i ��ܑ�����㼵�#O�2j��꧒1����'�ڢ�l�m�\/g�Kޗ����[LBj��'�h�k^1�"H�gF!H[=��f��6�4<��w�3�h��;�����o�K����n*���0�Wi�̓}|�)ΚXI`��JeL��a#iҀ�W�^fKx,�Q�'������^C@��6��}���~�҉ח�y��0��^4�M!b����^EUyZ���T4��"�pX�,�j��/s_L8H	ڸMfB�c巴b��#���Fb�w�u�Maˆ��rA[z�DK�N��/"1�ɫ�~e��l��j7��(pv��2߅��w��<ۜy�"��<py5r�nm;�����u��"�>��_a;�i=�3k�G�>1�甘�:�L�*�O��Yb�S/����t3���6/��|Z�0cAJ��'��Zu���ċ�ؠ��9DtK���*X��zʁC��^q�V�b��ڞ�Ej5�.RPk�o%;��/z��ѷ��۩
��X�����9?���S+��CY~){����ا�|����xu.o��<���c{o��nK����˽���g7�HQ�K���YW��������&�R��7����<�C��3[�L���J0�m*a[�����B��B�CӵS�2�:�״E�VbyB�Ɗ/Դ�OƲ�
�
�1m�k(@����]����c�e��B�E@������ڙ�Shl&�k	�w��̺M��'z��0?��v?�PPu�{I=t�ZH{�9�,j�d�d����vk8;p*�Y�����@�C�j�|�GbaE��XR�ƀr�?M�aa>C�zq�)9;`���Jk�N�*rO��(T� ��凎?��?���S�9}���pn���靏���	�,];W�������)J��a���{;}�w�o�S��##Q6n�#��ڻ���ᇵ@6���d=��oA){(R��cA����8s���k�$�T$;`l�v�i�Ů� L5n ��P� u��c�rs=�S�����}�]��v}�������ե`ꥍ����z��U�ɗ§Z�g9�.�������W���*v����W��3������<�������^���aK�E�yG�(�T�g5����+������e�6�R�	#�Ըf3&�c}�p�o-t�*'e7��+�)�)ՒV!�.�>��˜,S �w�ۡ����~���k슞`�"*M��9[/����������V��7�ć���JBi|�pG�&#��f��B�P�=q�o�P(�9�z�0S�1��5�I���dK��*��� ��J�!�}��,EM!z��O�\.Dg\��)^sD��\�4)(Y��]v���B;��u�Z�kŁ~�.+����i��nf� ��Y<�`�5��� ��v���U��T(W�%0���}�s�b.(��"�`��'-X��LױD~d��	heH�	p=/+�ϡj��ތ�P�M&w9f�v���(.I��j���;l�~z����I鑒}����b]oT�ism���6�����~�P��N���z�4;2�~�!��� �� .K�фp�ڎ����]�ؒ����t��>�B��F
���7���(����q�mv��۶�^M�}�����d��D�@gƵ.�k��
����2@D��&���N+IH'S�"a�8�U�A�ђ��XH��3V�o%&&i�[�p�:�1! 0��U��kt	E*�"
��;�������N�7�<�0�����6�LO$�q��ő
��{ۥ*�Z�+����55i��q��I?=���o�>��Kp/,�eWN3~{���P��2o���?��{4X��x(;���4:��$Ho>�|uS��?ʈ�?�w�'a�'�sd����(�X_*m�=�'�~��)���~τ���١�nh~�W���=�,;��Y>ݟ��5)2l���+�LP40���p��ݫ��6�^
%>�a�:[w����9n%���Ax�^�F*�S1����$���
_��j>���J}��������A�<gSg/�{bs]�Y\x�n䪝�
Sd,4H�V����f��M�O9JiOn��n�d�|�����}w�����
�� ��o6��c����Y(�x���f#���$��O�����6.��襮8���x�;�2)��D[��+�:�n]��u���i;Ѡd�8/�F��S�o�&|��!M8�~h<-��X��`����yl����`�n�{9�y�|`�Ԗz}f.���h��4T�A�R��4KpM���y$�%W-��
�^֧�3_�E����V�U�4�B���on���	��z�afWd��`|j�0k����@<i��?r+���x����c�%���A8L3?k�_W�{om�ޟ�^��a�`�Qv�Y�� �>X�Mm���>���B9l�b'{G�Hnd"و�\z	�o��_'�"�H:�7u	�ѝ���h���۴�i�B�>�	k�/����[�3�*��e�f�E�,x�ɠ���fJ<��lt�u"ajq�b�,sZ*�BQ�>s]]?�� ��jJͿ��=�@a�b��Z%A��/<�CR�)	R�ja-�,;�'��a�]�y��1�8:56z�I�/�t60vu1�!J�� ?@��f63]�rROJ��M,���ֲ`Yp�š�����$��"N�6�D
��Ԇ�i�P��W6Aa,�*��,ܟb����rD;�U�V�B���Z��KR������N�$��,l��^�C�%���I�p�"�>/ٶ���m��]��"s���/Os� 3_a"��\��S�|K��j!��"�x�2~�
nr�p���[�g+��q_�bR�<a"ɖ���^�;ʆ`ZjV[ɦP�o�oT}��^Fߴ$M�/�UѢ*P����^צ٦;ry&�K�Su��ˠ!Ƨ�*=]��m� ��c��eEŐOz���An�bjx�D��&䄅��p�N/��#|�S[�}�ٴ`gx07�92/C��U��`�-�̜��$И���%�}:>���,�^Lܠ� �_h�����:�"tC�� ?��=Fcj���i��Y^�a��k��R�|� ���U�D�4C�Š������RT�f)S���q��li*���W~���� K���6HJb7��G���*&��8���C�z��%�j$ac��j,RU��i���zh�+A��5�9:���v؆I̕lDx�������A��������d�~Ȱ�����P����LAC��	9���_�Z���ǲBś���`������",;���@݉��}uPT� Q��7d�&̚h�ks����ak��y�Dm
��C�����.�~�q�8��ǜ�u�����lM^]uE��'s�49�7'FnZ�\��A�y҂\"S��o��U»��}�3i���J��R@΢�z���N����4��c���ynm(��8g���^)l�:���:q�5�Ԑ1��Os�x����-�H�!cP��a=�c�S�:���h-�&B��@�$�6�{��N�B��H�]*��һn9�M�?	}aK1���� �������X��0���[n�\�)e�(�wG�Tj+SN�*KI|%.�4��$�f�ZĐ���w�Ez�ޑ{\�6%�WE$������Xv�܊�p��X��{s�ݫtG2o}Y�u�|w����b����5�]�!�����j"H�ͬ�������2�^�����p�p]��CV]���
�A/F{�$��Kqt�"��s��26B`��(ϡz���I���� �/�Z#l��b)>̎P��W����(��S���pÂ�����8A�B鸧����Ҁ{�Mh`�hA�Kuv���r���#����ѡfv�f��/O�Ԗ�����~��D�b��Úvx���
��HZ��2u]01L��i	���m���[o_��=��ޮ��sq�-NG�o�ى>��M�7^Hf�W����X		�,�py CFP+�{�t����C���_d4qi,4w��o�e�;�J����>ߤ�h@��f��~�?l)a�9]}�H�/5�8ӣ�p��9�IG�,�UP?��c�]�~�U%ꅯ]�_�AȂ�A{DG@���8
���o��Ŗ�2^���ιg��X\l��
S���%��x%!`�bTu�CYsNq�ZԔ�-�s�_,�K�O݁&�ޝ𥷟���kZ���EFӼ��[�$�:���g�0�-5K�*e^V�18S*����2�����{TZd�5��^�i�HR�*��`q��T<�Yz��=� �ܙ��9��e<�NT],Ԃ�~�3�<���}��7A�aAJZX6U���s�K�ψ�Y�7����9���rK ��#�_}�`�/��݌@	�d���
�We!���h����ۨ���j/���>�҈w�]��k�@  !-��!�'/l*��̚��W��d��5���u����p_�l��H1[�o)
'EFk/�ٿ���{r�l1��\W�u�H%��3�)R[��e?y�ӶnN잯H)&hO��l�o/��	|����\)��% �J�9B�����My7O�ߑ��q����[F��@��x��c�՟s��p��<Z�	�8����I	�G�f-uɊ+y��^��d��{�?	��e���I�VL�2/(��X^S�2Ɩ�68��[�\���k����� ��9[��/����p"m���Ù��HWG]$���2��q�i��l'bWI:ka�]��ǵR�ƺ�i��2L��^�	[Md�M��\{�<%����e״����p�lt�_R�,�F~�Y�K�9t��}3�_'{#�#m��:9�'��Н�ύ�=o�w���*e-�%�^�<7��T+#�o8�e(�N1�Bӣ*�K����N/'#&��� _Hj:��|j[ȑ��^8����� 𒯇nįM���x�KϤ,zX)M������"iɍmI�@�� (��f�J-���;'����oL�'���] ��z��JL5`3��V��<�!>lC>��!�JQn��Z�<�Ky�f��H��Uܦ�����D'�C��KU���DE�zô�������%�O��c�?�$5��}>��w�n/�j�;=l�����&��x�,�Gy�aGf.�aE��2��F�e-t@7�D�kz�E����|��L�����m'=��6����^��i�ly����ӤR�Dg����@>Jg�}�?x>��ݬ��з�į�8gHe��y�6<��5Q�F<�uc']�c�ܞHH�r��]���iQ���[W���Z|��V�x]>�yh �m��4�,�]hܤ2�i^C^�y�9&�ώ�Z���YRr�Ĩ��N�~v�U��bݐĭ�V]O�:n� ��J�_I�n�C��!�����Ž@|yaGN������@Ym8;�����3�N�̙���onuf:�m��a��!?W�I�eq_�]��oCQ33a�Wpz�y�(��Ʒ<��L5�46n�9��-n�vp�,��ܧ]�}�H�z�`B�z o\z�S1~�����g��	�����1�ض ���][mgK�<\���$�I	>~r).��(1�pF��˷�5������fS(!~�����`��"���1V��9/��r �^^/���S��>!��%��,vy���%���t.,�]�����pr��p��p����Y��s�Re��`-	����猕�L �$U�D/���´ףͳ�`��h$8/s��mU��H�j'��u�.,��|�����#( �,�;���2>���S�����:k78&���r6�&��9[n`qvݷC�8ا@2���5f��n�}��d~�t��j[������5�Yx��!!ݠu;�R�]�ԇ��5@z�
&�	)]m֋�z)G�0diN�m���':���B�&�����x���	ڦ^��P��m�Zq|(PL��;:�&��l��6�JzyI���MJ�?r{��]�X���,:͝�)�Jy�1u�����8���Tƨ6@���@�Mɷ�|EiF�]�X��K3�B����ҵA �!���V�*Fz�~]�0���OԪ�ޭH��$�%�1�?Ĭ�"t��DaJT`~FJDJ��A�[��$�'��du� 7q0��X\��=P���.�{g�7���T�((�	�����R?�9��xΌ?� X�:���J��vӪ�[79B��Upxn��T�;*�6�����ϴ�^y��.C�`@G���k���_�<ݍ�69�[n�Hy�(��p�C���I����7�_[JX���]*�/>8b��EPk�F}�e�g`^�v��N�3�9\����v�E��mT�NnZ�d�ɨ�Y�o�5`��\n~��b8&*�
�}G��U#\a��$Z�0do�=Y�/:�'�_Y�7�q��B���T>�w�%���G
~�sF�Y����5߉��1���EA��YQ[w �6�d>8K�?�'Ź��{�6�,%����� ���(y=��a'����n�pj�D�|�3*���T�+�i�4{F�HwX�WԎ�6&�{�\���l��1��}���ճCp�c�y�=�'>�ra�x;M�ޤ�$�+a��������!�D㗉����^��|~;���zc_&�0"
�E�j`|iOsx1�k;�mܽ�&Ǚ�a�f0�y6��I%)v�?���9J�����M�~D�@� �9����:�@θ��<��~��������ͻ��@����d f�z!��i����='U�"���`�~�l�`���uI,�bt�UZ�ܫ5n$(Í��b��a��}�pl��/����KU��`���!T�Jyd�1ϡ�t"�e��{�{���sM����M!�Z~�]\49��.�LM�����?0�4�@X���eI�ଖ��g~�J�z�����C{Њ�	�B|(|s۟��˲_�h�����N���-�m���_>�ϙ&B��������x]�3A�Vj%"���?I��N"�tq�V��A:��$�f�FF�^8�7B�V	���%(�P]�}j�W\�	^�_�q��a��;�A��U7��b0jɌi\���O��~��SH�_f@OA��@��rfL��CR�Ӳh�_`q��	��h �l㙾l�����W)r���$�ڿ@!����9=�V��j\ �e�sEġ�X�ɷT���['|�n�C�� �p��n��u�D�t&i��>�=�aE��d��`Ɏ�$�e;?=�pO��ȑ�|������Z��g�_I�@�xϻ
�х,�~Ǭ�����J���ݩ$����^��{�
4h;��NN,@X�/I������ ��׻�MJ3w��{�v��]�@T*Q���; �Y/k\���.ߩ>$�<�2̜*O]j=�|�i�x���N�p�	�7�f��K�o�G_ͪ)g�
15DXG%���h�"�5�=���F�?�Eh��U����*��������tT�`	����Ϋ��j���f)d��s2���ذZ���A�LW�~�HUn�dy��+��8�w��r�(�6�x{�뫺�7�]%�H��������ǂ��'�c��~E)\��-H������K֓�?�I��r{���9�%�a�#n�6��*\�cYv	�x�y��m�i��������8����[8P���Z
�-`X3b@h���\���<�ߩ�`���P�~�A��^��a�i˴�r�\�E����"�F���{����?�W�ù���ü(x`ٱ��ݿJ�Wg���@�k�������H�fȧ�	8iq~�a
n�8����Jl,�Z���w�A7f�� �(��N���=ߒ���U�e�S�bY^�C��a�g(��
U�	�����Is8��( �9�I/�l�݋!�1^�)]�t�(H���}��l�W�����CA�_%��y�����K�HG���/�7���TF�'ýR�֍KII���k�O��aƧr/��eC�ڜ���? �c�2�<�tv��uF^4�/H����I�lkɳ�M��~������#��T��1�UęP��q�wv%�,�������!B��Z5��|�u�W������IaF��V��Ŧ���oOz [��B���1�G�t�Fk�T-��,�W��l��
߉�a]J���YHUe4��cT�Dz�O!�U:_���R:?��#�w�"ǡwdriQ���O0��c��z��YGA��|�u�T�� �-fNB�w�j)��ų�|q����7�c�&"f���-�uY}a�܃�/��/��'	f�u�
6�/��A؟h�3g�T�;�}�t�w���cD���u������e�"3� �\G����=S�8ksQ�'$x����{����yEr_��K̝��c\༜NSF�|�aB�tE�m�gݰxX!������ߨ�m~C��R͕ZK\s�W��־��|�j#w��5�g9م�4Kya许[I�:�Zƙ�F�-`A�%��@�]+"��?��@�������-�&� r���A��z� yB�4�N�������ޘ��9�I�*X�V�.���z����::s�*[��nZ�)t]h�����jv�[N�Z)Lծ�Y��!!GD��u����4"�tm�y��n8�>]Nbt��4�
2��;�	;��T Y ��w��f�2��(�nEM�P�"�s!M��{�2p�x������<�I��mvr��!��:��W��8m9�>4!�J����
x�fG�ḹp��~��,��a�%|E�E�ƀ�$��r�{�:	�gP�a�0��x����0�[f�U��Nq��d�7��������Ǡ�@Ͼ&�Ư���;����`z��2��YxxP�b�q9P����dๅ���j7��P���?�Y1��K�����߀��z~�h��D��\e�-$��)6�1���@����mK�kg�
��Y��"�mn��Lf�L���m����,�eub�%ڦ�{��]�G�Ίn��x�J6���7�g�9ڎ��Ї�dw���o�/������*���6���
6��[���C�f�%軳����Uջr1-!6�j��i�^����+�D�j���4�Kщ�*|j4�bK���	��{�qk����Os�l�/�:���G '�PSh^�L�^��1�$(�=ݣ�Oz	�p,x�q�cEP|=�*2v+����� 7ѭ�c%͕o9Be.���-C��c������m�5�p�tK�X!��末k�������Ě�����D)��­uw���@��H��q ��gԎ T��;��a]Yjj�� �e�aT$g�8_�?����d"S�Ses��u�@L�O��8�	p��-Db����;#���w�v.�:Àl].�g��Ҭ�Ҁ۔%�d���|.tC�S�0ݙ������:����?XV��#�=l*r���d�v'�����P
6
Y,j�s�Y�9���`g��t���	>���^�W �0��UJI�l�_��a�U��b��_'�`~r�����t�l雑:O\���IJ�<z��J�2�C��KE!�� {��:zU��h���c۪�z�kp�ˌpz�X�a]QL"g멫h:����������X]�T8G�"/��C��,���m�_�!��k�X��L��p^�8���/�,�����3��n��$VN��gw{���z�;����`�uh�O�_N��LԚ��^z��:��$t��$����ՠ~i�|e��}E'�A�d2�~A���.�c��g�47=��3T�0�p��(��<�_���'`J��;�"��K�P�ʚ2��U�-Ȏ#q�Sb�PƮ�� 6�{�c�v���%��(@�>Л����O?����hO�N��k��,���gA'�W��_RnX�z��n� z�v��n�='q��Q�}QY�!� N��E��h�{l���5\t}
�_�ԫ:��@�Ҁm�Թ2�UH����@!���廜L#K�UX�X"��g���㨕��[[�X	�$�Y�ct�%�[%֥�g
�&��,2�fk���65�`�מ�_%�^�V/oȠ��E��#�e	!�A��xDx��L4�*��M��~��m�"|�*9������O�ڬ �d�4����V��t����OQm�7����OYh�[�Wm���N!JR��vF3?�������%QI����ʝ���U73�[J0��UĔ�ô�#� ���f.�VE���o8��Y��y��OW�"�a`�)��o�(0�����m���x��k���i��.^�m��_����K9Dv��_����*���M��ΟV�9ח#�0/,�s��ӭR �&��oB-�ΰ���2����O�?�� y>	�Zh?_!MiƵ1�)�X8YZ�7&IR(����x���%��WB�����m6s�p�_��X".J���*$�x�r���w j0ȶӹ*1uX��X�t̘`Ui:=!�A�G1��䁱in2�����5�#Y���R�� 	��V(d�j �B-��2nz��F&l�&�e�"ҕ��bݱ�1y;�*D��HoQ�+�Eٽ`;G�����:O��TW��iX��EAD�ҥ���N���ۭ�hDs�k�t�1̟����
�a�_�����`A��nG>'��@v]a������w�+es�j�n\��~<��ٷ����+�i��&�Z�H�&v�W&��Ռ�ۀ�P��4=�רӱ��M����ȡ[��MT�����*���@ng����o�������H�����+���K1�R���T���r�>���Һ.2`�h��f"�U{�#T��3������t�:u�3G�7�tð�=�q
!��>n3�p6N�%A*y��V�RN(���v%�k�Uj�����J�Q�V=�pW~��xe�s[q:6~Ke�]jr��j��U��uj��qnyL�7PMq������:�{���l5�A~J�wO�66q���C'ʃ� 1q^:�g��I��G4dT�G����1���-Z/d��xA���^��y�~v�b�H��Eg�-�P���!yY����^:������j$|�}����|�P%�T��8u�y.r�3��U�>^S��D�`�̡��Yc��E����e������@b*e'i�S����X ��1�24M��d�{�=�,5a�?��:����?�y�-qP~�K�<�S�Wʓ�M��l�NT���^��n�rü�m�2��.���3h
x� P}��q ��	=��K��)�<�F�ʂ����ڥ�����mPh^p��O5T�arf��}D����Z�Xف
Aq��9Z8J��W��c��G���T6�Q\���R4&Ů����ꄤ�I�:�(�LP_>1�Ԯ�����d���:�f��i�p��i7�W��+<%�K~|��Kپ�ULp�߀�
�7:rf�
%,�)�g$���� �,%5۬ҥ=��vbjy ��TB�#N�����y��m��J���������+���u"������j�<=����q��P�dȅ�Q�����$�2�q��'��ͻy��cY�Ym$���v�)��8#4��z[��n˟ϙ�"Y���{QC���\#��\��c�5�մ���
L�C΀]%:"�_��a2������fBn;-�u"k��ʛ��u�c�8�"̇;�`�sC�h�V�����7�OSEbCD�8r���Mg*d�P�U��3���{ͼ(�������
�Z8"�	��T����v)=�P�������{�	�z7'UM��P����T�Z0�j��}��=�tk�k�����X*�Y՝|D�V֎ۄr��ޓ�]ު�*��*l��B	���ga��Z� �Z�@Q���X��V�e�?w���Z4�{�r	�i@6i�n0��߾@��˧�4�8�c�S���g�Sn�Vf����;������F�G�� �����.���g,�Q|7w'<4n+����P�ȷRR`š���\8�J�N/3��\��W���,H�1E�V�j�a�N��l��))~�r����gDZJ�wp�O��t���^��&�l�3�#�!�C����Y;G��J�(0N+#4E|c������3�҇�[��eBS�o PL�4l��D�'	L�flf�f1��Zl�j����@����0� ���$t��X��tD�-��q�^��哓��2?�cǮ<����:�e��Zs�]0u��P�bDs�1
ʹ���\�G�$�R�	�p�h�� ��奩n�{곽�Y(ƌZm��ku޳	;��Y��D�a��� Q�(-��<��ݣr�����;�'�HF����S�	@KTm�ڎ���r('8zi�W�.�e����1$�V��5L�5�c����\m[���t{)�w����I*O�^_D�Z+U�p��@�*�g�'����.����t@�C�"rT�{��s_��Ņ�Os�F̗��	g\�.c��'��l>
��g��J5���V������X�Z15z��2���2o�v����� �^�!�h���*�dX;Le?;�J��gl��c���C�����$�Z�`f�3���"��2���E���]���
y&&��B@-��&�vnx̽���cl��x�5�'��{���Z������3��gҹ��{{�S���=�K"�i���k�+���v�x^/S>��#�cє�����Ã�gFZλ��I����Pc}V�A�.���P�]�&�f��[�+eQn�qU�N5�	��<ݧCqe��$�B���RlCF�_��n͙��н����#ħ�hoS{4��W(;��б,#�T-��7����"�����XQ�O"�������u0��i�\b����.��n�پw�n�P�7��T�r4��g$���Py�S���Hk��f��ʰ�GL��l�	�U�z��k!S��a�j��j5
�+ŷl�Ր(Z�t`Qa�a1��=��z�l����H�wRB���x�����%�ߍ�mA[�9�{�U��W�~Q�K;a���-Akx�m2��Wܼ�?l���g��!�5���_%�G��<���Eө>���@��s�-�F�|���-�s(�G�E3T��B�{�/]�
j�%�n��������W��@�d,d9���L��uIqJ��!�v/Ifx�^�dN��+��I`,C�o ���>M��_�U�ԡ�Pq��j�mϣ�>�Y�i�8�(B� ���/��U��A�h�br�'-���E�pup�`
�v�L���W���R2-w+���e��q���h��q�﷣��&���}
��mt�����7�e�7��$჎!._`��C�'SY�1e[�6�~N`�2h�.�,��A[���7L��|^��@15�ߐ{�R֗o��%e���qr�%�>aX�aY@�y���f��+�::�'���<۱�&e\\����pI��po�O����hG+B�G#���?ݼ��m}��1X�wv�9���D��a��B+9��]�y�n�ǃ�%�P���|}HHq�������Zn�|"	A��2�I���.����&ϳA��~�Ɉ�ŝ���@�Q��7��"߉T�� �E�W��ӶZ�f�pݦZ�3���ؘ<��
Dѳ�o���!WD�^�D,N���x�ӣ��������1*w1O~�{ٳ��/�LG��h���{�A �66���nK��� x�s�)T�h<Uˑ��4�� K|��R������@, CF*�,Qǰ���6�9�u�y2�h��ԍ.N͊g\ͅ(6^Mh1�6�v��æ�@"���q�N�D+!zm�A`�@˫=�R�e ]f��t=Y-*0�ކԚ�Lv9ڬv%~O?��C�1��� k�6J�X!8���Iؤ ������?���g',����à��~�f~դz��oI1�Z@Ǵ���^ǵB �\��M����@/��Ǧ�I���Yq�����P�Z3t�~no���-�8t��U<z袮����b����W��Ƅ[.��厾�n;���k�B�9ޝ�Ib�Og�ᬜ�x�N��t;D|��84Z�J����ȗ	���,#9�l�9A�꾩�'�)��97aj+�k��"`#���z���F>y�-� m�X����m��E4G�??ɽ����,��V��������c"��0�7SU� W��a>G~(�gPN�ų�K�?�:1��i��d�&{oRE��s���-\��U_ˆ5'd�Ʈs�L�Bb!���/L<�0��U��O���H��o\5|A9*��~��`��פ�ʁH����u��mC�*yF7���ޓ�!X�<�r5ruU9�W5��L�x�#�NC)w�(��M3	�6?[�ӊ�E���=��- fP3_n�-�w6�9���Ww�.ُkܠ���Y��?�����A'�V�#�{oʛtݕ\[�qE2P�C>9��Խ�!����I�g��=f�� �.�'͸�3�/���M���2r/��f�E��@9�/V���8JO�1�g'�+ +��~�J�fq��%o?l��شv3?����s�+���6��`&�b�yl�i���U7VU�'�Wa���r}����JJ�ƭ��V͖h�<�;Z�N�{�]���jy����]��\@�hN?��������D&�
E�\d����4��5��d��y����_�k��p�L�˰����粤92z�X&����J��ѱD��v��\wl�:H�����|�4�±���p��TP��̝4�8-[:��Px���A�a��ߕ�.��t�ק�--6%����fCO�� �\ʔf`'MM���u-W�+���W'<������X�Ĝ�Y��YU�2^�(i�klՍ
�d,�c��#�$�V��w�·1I	����ߓ'��
n�Y�z%��Ղ��0;�Ό1���@ÖЦ�m��j�s*����D]�E9�a�j�ký�W@e)���f����i��̅̽��U��0��i��}�{a�sOHv_��F�Q�4!����ę0�Rn�~��I�ڭ����c��겸���#��6�G�,���$���#}:eUm��M��
�*�W���`F�O�TQ�����h	����A��HT3���ސ�����cſ�ˢ���֟W��+:�%��p���Ɩd�;����i����+��6����˦�Wg}?~��9;�9mB�P����f�p1C& � ��<�L����R�"��6-E��
��V�	�`��Ɇ(��a_�����L����^��v8%��V��1���NYܽ��i�zV���m�x�j]Ffc�s�X���Uj�^X�pE��&j��ʰ4Qc����Fd��o��![Q��ͩ ����P�3�������|oC�l�=�I0ΰ*Fv.��.Js6��EN�,5�r�m)ћ-ږ܍��X��Bn���S�a��4�"=c1�g��~�z�ɐ�4>z�ȱ=��M�f�/W�K�W��Ʈ�6,����o�S�� �#oq���1.���a�?�)C��Ag���%q��i�6#|�^B������Z� �)qߜ�3띮iӣ$i��|��<D���U�d3�Fl�5.�i`C*������?9FD���u|�w�|�P��q ��E��&nUB��v�-����n2��I����dIﮨ���E�mc���?�b�eq���xw>�p�1�X#jV:U�FNT�Bn�#���n\�uF�z90U��ZgLCf��k0�=N�mp���7���B�l�r39@z[��g��>w;G��+��"�b�<{���@cS�}��-��=���J�9Y�D	�05�L��&�"�;��1�R��vk�K5�Ff~{��XlEsezi�5�� jJ
��s��'YP�ݾ�nq�>�k���,����kʤw�-"mbm.�卥�}͙zs��N���ps�/q��{�z�Zה�e��Jm���]%�����+��TlMȳ���*5+mK�|�I��]O-̮�,9����;9h7v�=�vF�C(�R����]��`f"���%�?��~����q�6����კ�W&v!���Wf����nG��r)E�؈Ԃ�5һg�h��Ԗ<�O�c��/S)���V����I|S,��	H[��w33�I(J�鸀����p����PH�_upV���J�H�"�a�e��XfzW�=��9=
iA�ϳ�l ,���{G����Ԅ ->�]�A덭3v��Ho`�Sԥ�=�)f^��;Ȥ�K��6*!��&"}e$���F8.��R��M�2p��R��1���rKOG����rL葩��(���&���/`�����>�q���S��I\�}�{���..v�[;j){�nl��lˇ���e-��	���ْ2�iX��8�Й� �Bn�p2�5�Mj���$t�}N�#F^s��<��y?��K��m��	M����:��E{����N�L�8��6�v���~�>E�������J���ߌu�#(XyX9�HJ-�NT 9s���H:q���[�Y?"��;�2pR
����7dб:�Dٍ|菊ψ$����p��QĿSda��)r��@�Y�r��F�����{���-1�L�@)DJw�s7��	�K�vOې��aG|zY�|��_�����C�<�"�u2�-������{��AY1b�R�ep�|=���ҳ�uGw.lj�h&'��7F� A���t�y�`�t�;�����]��3�޹>���7`�Ζ��Z�s&�'�rl�/���YE��*�a\�>[`V�Ѷ��R���P��8�ݹ�G�E���Ŀс%DN$������4͒��Ǌ���-e��/��P��F�SH9�k*z�^�?��j�d4PӢ�4NqLذeEP�9/*#$��3�����Q��_0KW��S����v�F%�F�n�"+m�f�h�;XK�ax�2�"�{$@���>E�FF��K}�-�a��� �<�����ǫ�+`�l�~��Y��G�(�Γ^�� �L�?��:��s��y�&̛ă���W7������Eo2'~���`ʫ[Ƭ<[+�������d���MI���Z��_I
룅U����k&@��Y���>�G橍�x�!��h��u�Ռ����@.n��%`53�L�6���1�}(a����Dɝ
%���	N�q����lEDL�>[?��{>�J�uiwP�4�`����Ξ,��?�Fގ��ĴRȯ'#jn��Do��PE�p=:B��������Ȇ��O<�Q�'Tc�nb��i��&\���T �m+�d�#Kwd	w,�/R>�f
\�耼��U������m)����Q�J=0=��i���S�BxY�	���+������(W3������;Md��@��J&}���|�YG눩���jt�6�5�@@�ɔ���HQ��~�aԝW�����3d�Ay4%٫����8��6��T�o�X}�[�HE��%hl��Y��{�~mӐ;�BzQ ]-!q0?��S�Cڡ1Q}y<o �J\�F' QW�i����C���L`��2����%k=����~r\�x�a�_�H- �+�%/2�]d�9���Xl��tkEX�0�Ĭ�I�ߦ�@1�q���q1��0!`,R����Qwo���-;�-�#�S�|��JW.,�P����_̎�6�dU�#X�W������<��f��h�nV[W�wX��<vv�QK��,�L��""AGI;�id��H����`���d"��:Y��b�_C��fqYd�U{������q_�T���G�*A���ռ4�h��K<>,��K���6�n-��p�V�(�������Y�+)8�U\&HO�����4z%PN8KNׇo6>��*<u���"K��4�,�:�1��D��t�d��i�W��S�%XP+"����V?,�j�S�6���գ��_N^O��9z�}�����ئ��URu�[q�Q�##�S�#�pਤ$B�^�9;�#D��`a�j|�V���|~$a�hP0�>��,&��pJ-��k�o-=w
���j��	�k���PHF���7ǘӛ.3V���R��^6 0
��3�ch�����P�	�;
d�����s������7�ԍ���c��gv�8Hk6�������Z���@�v���z�u�,�g��{ւ�-'���t�|�{�b�S��օa�Q>YlU�#��]����Z�Z�,Zw�������zr�#�%& �B��i��������R��e�x��B��}h	��ԭ;�����MGN7��c����%@������=���L���@�4|��P��v��b2�А�N
gO��#��� ��E��(}=�!�oԭ�P���0�g�K���c켂�1ֿ���,e�i�Ie�UǛ���Hg��n�>�}�����>��Aye
Av�/u��V�����T�<��Y�d��.d)�Ѿ��,M��-�a��e����� }��A��מiJ�����K:r�n(
;��37�M9�a%B��%�)�>��`"�^BQ�~������B�'�g�(+�	ܣ�Þ���tlK�P���ʽ���(����0pBU�ωv]X�����ٞ��]/��ܭ�H��8���xT��c�XF�t���(�l:��K&Dk6���������/���N�iq�6�|t<q^�8�%��uvq!��_��K��/K/������h�ѥRw�m��7 ۟�?�Ɇl���=�od*X$�v�˥��<s_��&�MKR���{�x"�y7� �|��K�_}%�"V��"uޛ`Y ��ZX��_ )����=��#� >��LF6��(S}z#D�� ����ˠ��0�������y��[i����*Q
<��T�@�S�x��_؉{�eud������vϗ�K��`�T��P���β1��)�+��F3 �+*_�*ɫ�Xu�y���`w�V(�ee�ͷ �q}��a����.sm�+���ۖ�9�bP���ݶ3k���<����>b��t`5ϩ�`� �w�3Y�ߋ��Z.	E�����#D���O�1�*�s�e[�������Ұ����n_�G{գ%;�3�Z���}��-��L�}a�I�Yv��k�kH1߻/���.��B~���C��RV�\����.��^�ռ	�ęa����f�N���*�}N�n�9���C�\�o�n��]]fur=X���)�o�dErW_���zVL��BR��W�Ie���#�X9��#t�w�,,��A��Lw�ܘ;b���f�u2|��a��~�|�Y��E/���x�Z��'e�|��R���x~4����Taq�ѯ}�%s��zlN��u���/\����gWФ](}�2�qW�*�*��a�ͺ��9�����[���N��NB���C�g�
�q�Ҩ�J�[�E,Y18>��X�θ��^�ղ�.����G\XSm��B��;�0��?e����@!��^��˾yRv�T��a=�d`Y�g�B��H}���i<�:�ʇʊu2��q�x��L�}z�1��6sڷ�=�~��K���_  ��<�FR_��0�#���+7;?,᰷��{��)׆���~D��;���S�V�H�"J����O�� ���v�уq5C�O���\ys��}.�
�$
�u�2������&�/��ƹ�YJ<3�֊�+�-����%�S��|�ʵK�D�z&?M0:0N�2��u2	���C���c�/.bY-�mk��^R���(�	�������뭃aS�._PZ��$�}-E���G��8]=GI�d��^X�?�F:}.�V�0A�,� �O���]���m�t�(B���չ^��ש&o���V+@o��t�\��p�����"˴��z`��}Qq>�����kW�!:G,�0f#�>�k�jX�P �zXɻ��^=��%� {���WLe�cI�>���*%߮���x¨��Tz�� �l�m��n`֩@�~x����D�w	A��I��D3�>�Ϟ|�c-��� �V1R[O����,�'��͡d+_�(j���bA�k:dÁ&+C,>��-[��2S�V�C��{���\�\��g��\b�D�(z;����r_��4J����&R���'��6fcO�o���i���F�:��zĴ5"���(�g�7�h�n�bpx�>�L��&�%�c�h:�L�L^���m<_�\�G ���}��i�v�r�T��.���J]XA��u�@�.׊��e��ݿ\�I�tlu�G�,7���=!��qZ�3����m)�=�W���?�6�Q�
}�e̘���];����r���n>Y�ɭ��F�x|�j���C{)mdqMuK���~T$�[�ĔA�ʍ�1ͭ#O�E<�<'l=܀O}�HLX��woM���.I g&0ip��:!-�ośC�>���)��?��$���=9�qn� ��5&� ��f�	�q�����J��}�d~n�%�[��A��g��6}V�q䆨:|d��w�w/o�_Lt0V��铨b��Ӭ6|��������x6���aȯ����>p�|a��L�s������\2��kvN����BC ��$�S2O�:���\/���ewׁ۷����Y�yv#��P�G�	�ӳ��]˿�ѿ��~��-t(�I�G_�'�F�pJ�I	?���3���,��TB��S�>�Ub| ç�(���:����6��|
ݑɦ�5r~�_���!a2ed�]Z`3`�(M�~3�wX\h�ĩv�������N���1�扠���������?dG����nL�4���_~~/&�}q��?�qT Z�ڹs�3$�&@U�׮@�C�ݠ�����1zj���H��XS�7���]�1�l���O�|��g�IK���[A!##�o �F/Й&%̶�Lw� ����$E�4����z|k��#e��v��8ߕ�����\p-?��{��Sf%�vQ����,:6vFM�*�$����x#�Y/-e��&h�^/��p��ݗ��l�W��~Z"��u]��I�����we��kR46��~�.� �K$�{�Aѽbav�/�E>;ܹ�w�Ue\M�W �;����Rj/N�_��8�8���xG%��Ą�ib���WR/*���+�k�#]A�&�L,c��Ywp��.��>��^ǘ�Ȉ�x	���	�ݒ9�E�:;a�n�bf�(�ڮ�pp sz��j\p�-{�c�h�x���m@0���K�JF ��>0� 1��a�Hp(���Ѡ������K��༈�S�}�<:�!b�\�>V��mHq�rP|*��ޔ�$:T�����L\�dQ���݂�,�w�^4|�=D�T��Z����jeJ[E~��� m�D�n;���i���G�f2�>�+�g?�������bpW/7���j�'UF>�1��S:����ўeG��sK_k�M*��x�'t$�(���4��E7��/K���w�{/ϯy2.UY�琍dי��ּז��^T�\1Oc� eD鏇d�<6��6R�%�=��aM�-Ї�6q�_(���.Y!<@C�hΐmj�S��gW�9�M��On�[t��dC<M5$/!�2G>Z�>���Q�.�"�wq���ڴf�@��m��ж�p�fC2F���T�+��8Slh`A�e����&�&u�d����$�Ea�	t���%rUX��8�z�����Õ�?��\!��w�A�>ɗ������e.�n!SN�7�� >8�4�@�����r�L���Li�j'En�S������k& }��I��H�_:h(g�2��S�5b��:VSN�
��Ej�/������=��>�TP�:n�B�3��A�ƀ��\�/-uW�����O��д�b�n>ğ}���.|�X=���@~l)�A���ǔ]���t�|x���u�XV:�v�W���C�)��F�?(���is��q�B(�5�<��?�����=��;U�Ea�כ�Y�\-M!p��iH���J��!�&C f���I����0l����87�[��*��(n����d1�Q>��A�5��B�`K��Fĉ�چ˪&y�����_��#���j��=7V��7���p��%�W*{���M����btM΀AB�#[
��]R.�hk߇�V�ٵ��]R6W�(SK��댕�g��,�u8T|<�ka�1��`჊���m�9����0��N�U�m�Ga��-L`_�2�x�i~�>�%�T>��@롙T�z�7�^�+�&��/�2�Ƭ��+��,���4� ��(�viC��g����f~ȋ>g���/��o�׷;��<�R��)!R��8�M�Wxol�.1�=�y���b��βِ���+F&D����B_Y��uK��Rŧ{�{B)>�	��a<![���ɉep)CqN+���JW�)�=��z��B�}|��z��Z�	�I"V�;��~�i���'����|��1��8��t:,a�:�R7,\fld�S1g��Y��`b��/��r�nＮ��'���|[S��bB����gHO5+�ߌ�Xcs��~��!�:�~��t�Y4�y|�*�]���)C뤷�f	�|��d'�G����jd���(��H��J?߮b�G���Pė4�^����l��"�����ʩHA�H�ƹ����@h���u�}��%<�u�ry���� Ǎ�FYW���Kһa��G��VJp����R;y��3s�'s�,��H� >�Q�K�/����1��:��j��j�f)��M�s{��I��D�@I��)$^�]���/=�`����A�rt񉇧ܼԄ�u�#��}b6b��0i�8�W!����C���B�Gp��ρ6��A/��m�H�.B����n��!�dq 0[��uP�L�l�ѱ�����ٮf��L?:g]H��L��s>UU���_�T���_�_��S��_'�~��1mM��a����x"��d/����m������j9��9�����IP�}ѫ�m�ob�s �ZK ��U��S��Ό��a��&r���)��Q���@rݨ�bg��U��hˆ����*L��j�X�\�<��>Me��@Ѡ��B@��N�tҜ3 ���#�\�l���	Q$�9:3���I�Jo�Mn�U�f^(O�H4<a�π�6���n.�r�ܨ��k��J;�0�����@iv�N ��	S�����B��b̍E:�ԩ)�������UQI���9�����j^B� ����64���/1)ð&i`|=w5�Y�
@�YDcȃ�>�sA���tWQ,w `ax�)�` Y�?ղ�u/X�VՑ�q�Ž/�v�W����/z��	�b$���Jȱ�2�7S^��q�w��"�u���u6���Ӕ���ҏ�c��H��.HX�س�.��h#��!`��uL�˰5x���J�{��������x|%�oCNMݺ�}�sq���	@�!��ʊ#8�>�v*��6.�p��#̼�|"���:��@��B/��-��+>�yt��EX6E�o
k�zG��e�9�7�7�\R�^H�p3<�!2I�K��A�>oI�@#Pa��m����Ƞh�F�9K|��֕$�9�C>�x��<Y���6�.�{f$���p�l������(��;��'S�{b���C��p/�$[�tĮ+Z%�o���a��r�����0���/G����K��%d��{/#��*0��%�Av�tb�����+5ʺb�5��6P����b>�g����軿5�]#�?�{!X��)���m�6��_�?L�=��^���dB����#S:�.3ف�Q�ѡD�˾g�j��Ή4��5`-kA��%��,�P�t�/4��d���W���7�f4ՠ��oڶeM�t��J�^>S�Y�F�2�˴j"�;z���"~�-�"[�G
�5�Q�|��(�~\t$я�E��K/0�R� Lu�K�T	��n�d���ى��2�S�����C�4��ٽt�t�:X50��й�3�*�N��Al f/�@aX핝x����|�����U@O�H�U��(:���>)u2D5rp����+s���L�#�6�]���N�Wt��8@�{��Z�r����M +�X�?�l�Q���k����DT�0H�f�<\�v���f!/�C5�1��#�95���|�����5���
Alq�<9�\�$�"�̻F#5B�FUI�<8nϏ�o3W��0�A*�ڧ2:�~��}.�BE[*��zЈ�!���*z?��E��{~]QG �;�����5�hL?��ɀ�%�xT�Z"������	��U�5�@9���ȯ����y��B�F�>��U�l3 P,ACH��z�6�""��r�\�]�����_���I%������c�R?� 9���
𨇲
�O�z��i�H���C_#$��D����~}T"IK�}J^��5)��j'd��c��dr����C������84��=5�U|a�� ��&)r�OI�Ho��֧MC������W��R$�����_��� �F���['��eN�L��B^��ݣ�3����C�zy�"SV�Ы�b��,�-��<�T��}�;�:�$ބ)3�A�'�����.	E+����M|�?�{D��3�\;fcf�}�`,�an�g#��9��ԫׅ�.���EA:��{���@�;2��v4v?)���<�"nߩ��R-EO�C.�IRbqF�f�"R�.�.�٪�Z[}gX`��\�O��u�����!����U�L�c("YF5,���v��[IZ�T+A��Y��y����NO�`����ϑ���C�V�2S���x\`E�WӨ�籘a���nV���C�6=��z�E�cs�mJ�&�5�m��������*�!�{ΆNf��G
�����{'nL�2��_,9.P7�~�=r�ҝ��I���4ݙ��!�b�߄���҂&v��!5��SJ�x�y��v]��O���O}t+��E�j�p�ȕ�j����L�peSwNy,!>�P�G7\ut�6� �OQ~��4��VD���Z\�]�'1�}��8�.���M����W��*�"���(�qL��$Ѐuj��	K��D�;7�u��B~����eG`�G+n��jΠ��q��൳���Ǭ}b�G:R�����K{��HQ�/ͦI�S`�;!Ȏ�kM�g�U=J�3��l(E��1�̮�>��:ڜU���u'G��Ek^9n����x�z��l����F��m	-B��rl���,�����J�rD]�`s�B&��a܉1���C�P��"�x��J����u^�뾬� C$�J_�-^P���s*���yʙ��<�T~`�oV��9	�G�`~�
���RמO��	�+�)�Ր�n�)�FA��	�n�s 9x��ն�5s�t�-N�kN�$�Rsq.A}���������ꎿ����~�����O�~���#F����g�������(��c�`�.�:�d�-N�RsGw��OOw��mm*_�� \����{�<}��-� 57"�;��sC��S���y4k��X������ �?��~1o`?��.� S���ul�w�h*_� ���>�*�S%����;�xu��)b�I� 7�� \xx�����oX*zQ�慩�k��z����?��0�mS.0������k�ϟ�X^)-�d9��&ʻQT�,�eވ_��������tz��_ PGs�����?�������~T�5Č���Ms@<�a#"������?2�t�RqI��N����N�_�s��a�76��pJl����=ۈ���f8ԾL��1��mI�Ď��ޘBY;�N��?F�+���Κ)y��?���[�L����!��`��1lȎ��*��l��1�y��=�PpoLK!���+��7]~β���h�A���^���rUo��+8oP�N@鍊9ɫ�±k�^-��_�6H��wF>�g~�M0�h�����@ka��W�?�h�Z�&��q��'?"�'s��xq��S���oo����NM�D6#$����/ҪÍ]I�X��/��'Ⱦ`a+gf�r��[���O(C�$�0�t�8��P��́��Y6B�=d+��J�� ���\£i,��Z����_@<_w��nA����_۬��QC�am@N�#t�k򔜻�$�]%ֻ�)K�L�U�/0R�I��Q���n���
��9y��B�᠁��eG0M�3�	�`_��Ɋq�b��s?��`����g�a>m9��c%���A��,�<+��� 9��s�s9��y`���(0O��;��M��l���� �S�G�B�f�E��8f�6��T�v���E$[;l\��q���2M��a�I����sgh�6�9YG�;+B<W0���f�&;Y�ґ^~�����ܶ�v�?�L�QW���3�݂�u�ʫ�{r����P*I�0X��g�����d;*��/v�4ia�m�Tg�_/s�da����(wg�at�*� �7A�M��'�7��7���w����ҁ۱*%��f �*q~H��0'�,���-���J�C����!�C�����X�yzK�����+�1s��Ôi#��5
rg�>�>��nܔkI�I�����v���ʮv\js��9�&hA�Id|���˥�%�.��9���^��Y�a!�X����k����N�����xB��hક���`���ܔ� ��[�H���D�֎�F�����,>M�w5_�f���j�p�����z'B�Hc��������f�J���t�{�q(6��d�{z�V�P�q�ol?8�B�S���8X��XS7�SC��@�y}Of�I��W�_AR�OG��醋0��6�i �!/�c:#uK+|�,`�aR�lT�bN�"�!V���CX{��_XM�mG�,x���d�Z��CA�;�Ӕ��34���S��k "
_:0`]a�A�O�|��xɮ�R����K��kdm��\M�y���,"�*g�f�R���A$b�e���`VȚ�[�N�ya�Z�A��e�GI-2Ez�U�s�xo�ta�����VZ��ʀ�i�lhl֧Q�B�K��%pؔ��Mm�̡oN{�o�҉!��	lG����J5�D��|�/�62;���j|��M�Mi���ZV&�}���F�+pc,��DgY���?lA:�	bM	rJn��P��t,1���s�Y�W�;w%���'e�w����$bb��� �-��P�T�*]�hR
�r
�=/y���.�����*��pjB@-`�q�����37��]�l�t��$-���
_]XO���:ʆ�cA]b�Ueh�mw7�p��W+A%�y�r��ևv���3�g������"����r���Umb��-O�.	��:�o&�o�X�����m�zWۤ���ǆ�v�8ʰ��`�Y㭝����=�Gғ��(�A�y��q�蘟�`�/���B������Q���t��8t4sj�m�����ߕ�s���-�Y�pq�����$��1�2�����t��1�W��n�7�	h�ÕF�ޒJ,�k��4*j��?�$���}��E�F�\��hDq�:����:Ո*�)�c-�_Ǡ��<QQ��*g�ip�X^�U�Ol�͜t�b�B@���9 �AC�#�iXW-;3cD���I�.V��EC�'.P�E,�)����Uű��
�w��8�5�Di���#4�{�'�N��� Uɓ��Mݽ���E�O5D����Nf���{b ���z=�˄C�֧�����)�o?����*{DDپ ��Q	oĦLnŠ�� �|g�JB;���n�n�>�I��7�|�S�����B�H��B�.&��_���`~}���Po����9)_uΞp�ԩ
b�b/�Fdr��`+�cЗ�ӂO��.��%	rgt�ET'��&� i��䕾����F���qF�~�E�(��h��=�l��(�@�e�ɰ�s���T���UbS�]@��l���)ziV,��9�wP��1��C���X.sv�ll?�m��uO륮*r52��4Ss�]Gy��b��gw��V��g�����[�һ���q'j�h�|B����Յ����tli�b�,��6e�Ճxd��93hQ�وʆۜ|l�6����AK;��fy-�E��_TWihu���|u�Z!�<�=�p�K��-@�~S�ϳ>�� !8�4��W�_�p�@&�7�_їvHH���C(g�!?D���s�Tz<���g�?üꉲqE]����j��[�K���9���J��q�=�W�=�Y���1�����m��e�S���n��40��HЍF���ɞ�T�?�`�د�)����dN��U��'�x�86m2��Tﳢ{�Ո���2pQ�|�*�n�Ju�;����������2ʄ�L�����]���ǒ�{*^��~�h)Q�v��(k]^]oג�"e�P�\�a��y��"sB�s��/q:S\�����`�2r����n�IqP\?����^��'�\���s����2�i����f0y#�GsC�I�PLl�?���)�Bب�
���N��΂�w��Ô�/�'z��C��,v�9 �S��S��3fI�Ê�b����uN���;!���dꙇ�&�ј
l�K��v��%'�Wc9�k⣚�x<�0�%<ͪ�?��9-R�L��w�+��z�M*Tk(��1�연�Q��$��`�F����֯�U3ӓc(Io�T�+�j9^��:9Ẏ:�\���X�P��a{��EŊ�5� Loz7>����v��WF��B��^��$��ɾX�WY>NhW50����KH�qZ2tՔ���o����k��+m�
}F��\��EY���x6�A����v��r�s-�5�8^Z�ĢP������ j�M��`0�ψݲ!��d>�D�$S�u\)�����J���n:��o�̙�^ݱI�d����~ˡ�Cu�)N!�����Kk0@�Yh���.��L��� ��tI�ܞ�[���y�Q�6$.�Ƅ9�]���b�0W�w7z�SV!��)�*�U#��M�V�6=HH�:�['N����[0�؅@	�h��P��:��au�p�/f�QSj㨏%;S,�6��W7��@�	w!1.3��-EQ�`��<w����A"�F����\$fڶ��b9P:1�Rf1�nr~ܦD�#,������)�=%-��5��K��SG !�{�r�:�4[�9X��g:��ƻ	_|�\KH��X�J HƮJ_���[v�&[�;�m�@_8�(�n���)J
?�ق��8��5p.xkZri�ͤU�d �e1ݓ4O�d����i�~Z� & sG�f�HY��U�uvk0�W������;ё�sI������"Ыsd@DB�R�a��X�����|��=`��^`�BxĐ�u�W]}eǞ�e�����j���6��\�G������,np�r���w�T�#��G9�ҭ��}�TR�҅��>�DT�Wz<׏Pːb��͟A:���ޒ���W//Rd�D��r��v�S<m�\��gC\�b�tU����[�G籑���ؔ��d�bs��8q'T�G��D-�/� u=4}�#��T�y�O�S�!S��pA������pV�8�� ��͞�Z3���$�s%/GL�bfX�6����&�ԃ�TR��k��W�g]���*�4�w���p��}4z�B��W0-�K}"?��
�z�R ;~�&�\w����Տ���I��G��\/R�6�<�,/N���~	� iw�cwY�A5�gˁ>D�0_�L�m�>��fn���(�3M#H��uo�֘��Y	r4"-%P��"X~�a����P"yq��O*�ZTO��x�B�`���?m�Ź@֔z��XK��қصU���3�Vea���ʻ�?��g�GǦ�M���
o�-�Iџz '��ϭ&�{�jDCh�'��J�u9o8T�N/ې�"4�܋��nwE�x��Q�.�T�־h���Z9b o����QY���V�M��*��v9r:Qn�d�;���^�h���F��'O��e�-w��>Ŗm֮8��.Oӽ���s�{����|A���T�}<_���y0�o��-E=wN!��?o���y�"���ۇ&$/9���[�"(,h���H!2�|�ij�e�_$p�(i3�An���H����4����o_[��C;?ƌ^3�ZN�ctqz	Q�9L�nk}�����r�(�HW����gB{�+*�oZ�kH�Cr�L�⨙��'��8z	���HM��G{�$4��iЉ�:�@�� ��w���j�����߿�F�ɶ�����p��Հ;y����������� -�����H���4=��D��TTv�{F`����pt�]g��L�	�<A%s o�@>vЌ���6f���s��U��/�߬��Ή���Y�_�OP�;r�����;�
�	��]��V�2�2�-�S^�1�@�>W G�V��7|��_��3��@��`��n,��K�����$@�?$�`?���4(C5\r��+D{�Q�RV�r�mXN���	��'��L�<1Pɩ+㰓.M��O��&�2
�Q�]0g�M���-����y^�@�6 ����Z��I�9��'��t��u���cy����;`q�+�Ѥ_����V�=8����tčJ��	����8=�ݑH��_�o�/�ٹ}���,MN��EAF��2-z��j!������(t�Η�fd:K�w|v��I��ύ_�sB�	a�i�\�c�!������G0�i��"H�[���hq졆�H��L�5��i��`K
�_a�c��r!�Кg�9h�'���΄�j�D������|��v����u$_RUМB�
!���6N�d�T��n=��Z0�����e�Tx�{�@�~2�[��CR��ӝ�!`��+MQ��ALbLH���1v��>ِ~W�d�IBr�����+������?HMu&e�o2�_��F*Z�_��YpS�17�F���#����BԏG"���F ���\q",zt�F��f�&c�\O9g����w1B�j~Y cP�L�����bY�#!�wg����d��l.���G�4����F��Q�EiK��}�tA)�Wt7����� 4���ݼ���W�YwN"�TN������]q�B�`�#���D��H���t�r
�lS/��0�[�>�,As��!���d�H��v1Ũˬ�{���k���Ο�h��wc�ҭUhw�anD��W����6ewP�7;B�
*j=QᒺD�8��Y8�$�Xa�k@fik���8�״��N�/�֚c�;��O�[Ę�����L���K��cNPu�0�}y>��KQ����=j�/^{E�^�P	��ن�8���i���n�����`v�c�XB����ah���8Ún��Sstb������3��9}wUSAvF]>B;E(A:�� M�Bv��lR��8iZ~>	p���}�E�ؐ<����JB�ꃜg�w]��[@u�s�XhR`[
�a�VN�3�Ш�N��#Y1ٰ%i��� x˧�q�0穌.��u���$��&�-����1/��pi��L@�>~��S�n_�y����K���s�(G��ip<�lA4AiM_���xY5�d����H`Pc���:���Q�9����dD�N"zӐy$%D)^w3�U�&�����c{�/���)��	@2b-j[�����v&Z��j[��[!P�<�M|����-��Hu�ْ�d���l�K�=RU��3��h������*v�n��4֥мd�����æ)�}II&H#����SS�φ�Ƚ��fy8p�7����/AH.��e�q�lX�3�!t������qQ�,�+t�k���[�{����x�4ٖ��� �Q����˶�!KqC-��q���t���@ly���Y,1�n��t%'����"���l�jW���
0-�HIǖ9n6+�:hM���1)�²3/�;�4&�	��U�y�Y�i��.�W.ד� ]��� A�v����L�ęґ㪯B�0�������qU����et\|�/o!.��/��s�`E}R�=�RqYᢐhQ�F����+���B������JG� P�������N[��=	Q,�4�A�9�tYF7�яఽ�� �����|W�����Z;�U�gd�oC���*<�}��3,���昲}I�U7@3��$h�l���a�ٚ�@aa���%����}�.>~T��o79�/��"�`b&򡶸u���y ��0��CR%���1������:|�C��0K�YIߠ���qON��4X�:K	x���w�p��]�={Ӽ%B;?�����1�-�����Z�1V��c71xGϥ̥����J쿊Ôj����`v�"��{V�7V= �s %�۹V��b���c����� 4X�|i�e`������s�(���� ��(�f� l�0�&ĸ�aD[�g�-Y5 �1Mhl\6Y����3̟'I�u��y��uU�V����'�i�X�;�vZ�a҄H�ɬ��C,+��d���J��c:����|��z�R[�^V���#0b��7!-u��69�!\��:�W��5��KT6���Y>S1g5LwQ�a��͌w��Ax�˪�DK�o
�޽yq��&-��?wH}fc㧜+�����*)�I
 ���E�*��B�A�Jdo!�k������O*�Bq���e����Ե��I�d�a��Њ��6w�G�_&[QR;�@���m�`�|�RD���$�Iq�%t�Sщ*Jx3�|ZFLN�l�i�������@3.QV�n�E2=⿔v�7wl��OD Ņ+�r�o�#���(�K��CX�O ʩ�C_z��D�f �9�}�dj���<��N�W�E}�Nr�G�����LE���_p-� <�ʽ�#���"x�K��F�S4��Z��tʭ%J=^�:��*�"{�r�f���>Z�sS�`6W#�Wj��XT�[�������_�_C�V�8��DB2�RwHe�������?߾B��m��ލW˫�XK<��P�	���Ul�>2�bM���W:�r_�{l8�Y�4� ,���*)(��th&�*��tӸ��용St"�p[R)�,�rC������-8Q��Y�)4�۔�b��#�?8�^�J[B�=;�86B%���s7�����lL�98�Qȉ��S�?O,E��qى�������>�<��)n�QB+dN����-l��<��$�g+n���T��� [�K��bb���3���Wl�t⋅��h�<e?�Ӳ���tK�.���fx���b@q��d�a�n�Lo2�c������Vqu���4�'�K�y`���Ka��s���(�w������$��ѱ�1�n}��nd��t��i2��%��^�{�j����-920��1�5�y���Oa�����}����Q�]YFH�x�s��)�ueI,����~=�)c���y�0�E&j�{!v<����pap{(UJzfF8��^�� ��I�}fG��� ���mVwd���T~��١��^�d�b���#*�Bʄ1���!�3-� p߾͸�a!j�B��]N���<x��!�
O�����#bH��uCzʪkS�FD�S���j ���ݏ���v�Oپ�?E=@۝Q��xQ��N�#|Y�(!�fG~��喙T��>���c��͚>2g��ֲS*V���; ~��sO�-	Ҥ�5���2�`ޝ���~�s�� �"%��>�p���͞ܪ!��d�O�r���IO��v\�QNW�d@D�Og�*y[�1�/�XAI�e4���r��$�i@Y�]0��;�z�n�B�� �"2�s�i��g���P���x����$xù�(������"y���I��#{�߹3v��P��4�`&�F���$	����5��,J�Y5�Y$.WA���W�)>�U�j�6I��y���dr��;�@�}��Y�+�������:�E�s���D[�0�={�e��q& ��D�����蟦xIW/����k�6E}�5�4�I���Nͻ�E���e���p��浯�E<�pV6G�g*�[�^7��`��D��Wpp�'�7��V������gHĝ�DT�e�	�
p<��'U�� ~�ߚ����r��3(����jŽ;��B!�y;!h�@�9n���K�<�M^ࠂ+w#gP��E����ڑ�x,�d�dn[�	�$ 髧�	�ǝ��8_2] �f�U뜒���W�.٭�Rz&	>�ǟ�J��<N�{}�ªЫ�%��Wk��J�Q�.�hы?�E�(]j rV��Ѩ�AS*��h����vHt�k T��6^��QD��l��<'?�j�h�)�����?�ܙ=G(��b;=&C��v���շ{���ߤɞ{mT�ȶ�I���*OU���tKȐ�3{�Ip*��0K�6UsV��ٷԛ]�>S�*w�=�WՔ�@�`˸hi��w\X7�;�!B(�I涁��Vy�k1bv���y��)����+:~69�)K��Lh��ka݉� ��+�!��W�S#H���\�&�\�o��۵�{�p�(���MT_����~�'g+]���S�©��o�SV
z�菦�l�F�)�E�5�݃��{]��[j�UF�4^_W �HϽ�=��3��*f�Q��oً�'g�,t�A�&�9y�o^��%_�{�Cn3�#L�?�
Z;��1D%Z=��Hn���e�OR�O1��k> ��R8*_�6ov	�xB�ۂ���M���t�
U����M����SRC�=�(���M�Ag"e{;���H?Ї����wHǱ���=����
UHB��8���x�x��U%Z�-�i�ݧ�Ed`
�m�k�J�v��D3Bʅ��qU�*:��� VD�J�t�-����k04����S�Q=S���Ay�>�����ǾӡbZ/ixV[;�CKG��K�Y�XkV�e#�],�'�������1���}.���{d�����Rf����7^�̣]@�.�\�Eʞ���2qζ��1��OFv��_r�&�ts3�Z	��Yu^�[v���>���esb+v����-����я���8TQ�R���p+�X�Kcٞ���Z����ij��z��ef�Ԍ��j���Mꂘ�g���:�V+�DRȡ��C
[;���)�Œ� t
FD�_e�X>xr%��e�幛�,��������#c��F�H����	�g*Ik}�7��P-!%z��Q>b��M�"�\Y.����\G>��˟�������7���2-����h����R�[��"��Qw���l�܂���Z�9�o柺�XQgʳk��&���ηJNc8�	�@��q��Yh��\�Y��F������m�*�� Mm��� ��D�'S\n�h��/d䨌K�f^��Y$�&�Ǵل���2X�X?���R��;Ү���H%9����T��܂�������yP�|H��[��_��$/䃅�Dj�b���A�ȑ��ʝ�VP���r�V�a���s6�0�BB�6cd'B��!����G12�G�u��8FYx=�~���Bn
�g�t��������hs�6�<�0�%��Ң��Db�Тxd�Mڜ�ơ�֖O��ҝr�nw;S��f:Ȯ��0 lDź�<�K��e>�ce�Viqa!w� B��^�W��3}�U�@��W�x��s���y�x��9�V�L>�.�g�͇O��;y��'�N�D�aÛ�5o.|��)���1+�$����9��r��k�G1"�<P�-�g�U#����@J�[]mX����MV�8�W�!� �Ŷ� #0��-؉+�)P�-U�y�7AE�s1 qs�����'�F��3�I���`���Iڄ�GeLK���vǴ�4x�0� !�R	r.��ާ7��h��2zWq

��]pwA��`�,��������X'��L�1������G�i-"sI{��%|�� e���]��{�I	�@�Z~V��|F����e�t1蹒��ô�M�T����Fe�@��
N����8�=k�O�Zm���koC{2�J��X4,��d}�t�0 �A�ߵ�6k^�ѭ�n!��|1��A�ߒ&oc:�ao��on���!���R1m����t�Ul��G[k���iQ	��]��t�]J5���O��iG>Ɨˉ��x�Gf7v��^"���LX,���,�m�i��E��p��տ���b�B���l�*���d-*�!�,(��H�%�F£�,=�Zz�'<�l�����l��񙂁�
!���-��wc:��HT'>v����%S[�Q���F�����d�ޏ��ia!��'�(ycpqRa �~*P�I��o���J�4{��ɺE`On��y&e|f���+��b?iuS{��sa�!U������G�j���-V�n�yq%�G0�HT�M�����͵�b�g�k��f��	W��[���S��}��l��_�܏ %4�V�`f��G�PytcYE�u�"�2��1���H*��������c	n���"R��s��'��
'�v�Y��XU���jE<L��aה�U���֭�.xj-�6� ��_|��]���_�$7�s�d&�����Y�I~c��'��H�Z��N;�	�+�d������;O���)�b���l"��I���&�ࡷ˟�V+�6{�Mt��r-LQ����WF��+`k*/�����dǎf�g��#�(�k�'d��2����9�0�7�B��1��p���M{��߲=�u����}�g/mB���7-�Ōf<;�p��DiM�;i��Oc����j��<�x^"s \
������o��>P��4����U���,�����u%�ֽu��óp#�ٰ[o�Q��vS�F��Mv㞑A�Y$R����a+nk/t�S�ֳ��R����<��+J#�� ��x�)3����-�`~@���$�#��R})W���]srn�gb�����%��2��_��0L)��֏#�ӧ�4Xl�4���5���N*:�*��8G��T�j8p���[��[U�u)p���.�����l9�z�*t�U��d��!3�;Y���sb��6����9 5p��#�{(i��h0�X���x)�Ŭ���@��L*zZ@����I|��0�[]��9y��&~(�mþb�z�@��Ƹ(�A��N;g{��8`�]���w?�����vt��@*��ȇ����{�ɲ9ع�	��S��La��s��	h�x�ג�ȼ]��$g���VF�(^BJ�>"��F^�����K����>�����pQ2P�@Ù���O7�'�; ����轐�j��x7�����1�V���e�yd�pn����02䋙$���#�Z�dh߂�f�?^�+\�
{S ��`��{��ƣ"�#�S0Tc0K"3�I���+�<��C�Q`G�:E���W�u��f��.R��ɋ �t�t(����0$h3�YՋ�*����[#�B���g��U۴��*��+���N�U_p�Ki��b׵[&v�&�6K�^��e
�;5Yv�4��d�DhO�(��O�����c=�!e��*��mȋ�^�"|vV��h!G ^�*҄@̄�T�Q_5
�A�mAs�S���:�/�J�X��yPD���=c�cЛ�d=���V[��pGI����V���p00��h+�I�.I�N�e���<�y]q�������������B�k��[΃Iҁ���<�2�^��4���ސ�����.$Ľ$�^pѢ뇿��(;y� ������tO�����^���g��9yŴ����P�	�r��XM�3RNo0�h*h㕨y���Z\�.sa���,R?q?�^eB�Zx�ra��\.�[�?�ܨC�/0�0<0iQ�_���^`6!6��d�|�/�j�nu�R4���W�\p ��'�L[�B��E�9����vv҇.��[�����u�U����|��r����R����ռ�O��QnN!:��Jf���'.�DE�r��T����Ett�?JCڜ.�G�'�LM�tm/��iK�Wt���j��/�nw��)�����nE���^jC���zkO��~)Τ3P�v�����r=�,|鑆�K�aYX�blJ33O�}W9��o��f�d��Me����~-�����J�j�.����r>��Җ��t��� �m�ՊTe0���k�D���*ԋ?i��>sU�M�`�0�~�s���Z��i{�ŷy>�pv�v\�e��	]P����m�t���t�?�@N ��
��}$	�V|��ߡ���T�b)Y�=��v�(��%5j��W �Kث�?0�Y�B"lQ` N�#q�|���ybĥ��a8@5�[���Y^�<�U�Vi7�oj�z��)��O�X}'���-�iWj���:��s�����Ca����ۓܕ�w�G��TC�BӮ)���#��`���:��BL�����Di#�]���6 8��m�]�P���[��؀7bBx�?Ȳ��zQ�
3:;[T���:R�f=$��(�w��?��qV�������I��wAʈ�2����i J��r�fZY��������/K%���I+^�
��Hu��=��i��wT�s��Q��zg5C`�[>dm��k�+?�B���y�W���?��t˓�q��`O�Y���������NN�?��]��&��3�8'��9��zSTS报!�����ͣu�"��+������BA�U�e��!�;���\m���o��P�̀�:��3�y48=t5<Հ�%D�7�r�����!�c1��j�(�moPE�ƪ���-rSyI�<N#�D�:���� >��2�	��Ûxb���c��?�@�f^-���QTB�'��(<;�9�+R��}�G.1���ޅ٩��C@�&�E�%�UVi-�T	��W�,�f����$��d��T���s.s(��q��ɤ��� ƿ���)Ni�y���E��a��K8yKV�.���l&�3��Ɏ0�^��.���S���b��p{��9��`K9g��l_$��>N��Yn������I(�Q8�������aA��sPr���H���4�g*v}���C������	��)�l���y��%W�c��װ��coz�I�_�ܙ�F���Qg���(�3����[���Uo����,�%=�5,�s�|g~lyg�����ȹ"IĶի��^=�u�,�	�%nH�ݔ+��E���T-�"g�xs���琯q0�������fO�f�6ǹ�����>Ȇ*�e#��@�V�\�`E�/�u`ڼ�Nb]c��+y�yUMv,pt��M�;T4�[B��7�4"?��;�ȁE�Z�X��7��6�8k�{��<nj���D��|#՝j䩾�[r��j�W����Y�89�"�U�
mOx47
hT�8��d���� K�_�Q�v�T��&��eA�\�����Tg���i�/���d/ʅ�/�?�FG�z4v`�ص��GD�����"�#-�7qy2/����JN�M| �J��3��;�]4�˽2fJ��k-n��0��"6W�Pf�0�ߍu���C�ܽ�X�$�9�K ����̹ ��P��L�":���p��f���0�ӦT�M�j�DǤq	��ez'����Ɵ��%�C�n[��#��ב�R��3��?�P��4%/�	i��-�7@߼$����Z��WfΕC��7+%�Z٪�� ҳ9ͻ�k�x���!�Q�a᥸�0�L�>���"�7>������v��9�ڪ��lpP�c��$	t�!z+��k4oi��LPED��W�v[�^Z~�`����V�l3im	���~��l C/ҟ���)J�܋�Z�+��� �ۧ����D!8ho��*��ɯo���M�(޷��S�j�ԣ��b�� 4�Q{��r>��q��&��M�a����������~�����x�4�:y���o�$����������FB~6}�G_�'/^���?8���C�c�Sʀ��S?wBN^9z�uUC�՞���V<��P��=���I���P�M_��BT�}�4���52�����3�k�eu��w�
�I�p���B���	y��@�	9��x6ƀ���RX�e�Dx��s�cc
�b�)���q������6~'$(�=�^I��*om��j��sJ�kWX8Ϸ������('�.�nd��|. ��?���|�s?�d���,:I�Q�X�Z0�_"Ǵ`fE����8F<�p�}��Dy���y"To�9Um\#ȠS�I2ڻ�OcyE������Q�~�#��1?�l?�i�Gߘ͘`����5��w={����)�f8r���;�˱R|����D/��>�]0?d�����ө. �C ���.�+L��Qa��F�W��v(Z�\8�,��&��1
e���(5nXT�vQ�;鱄�,z&�no.W�ٮ�Qj�ģ�0��|\��#|���E�p��-�D�Ԯ%dE~!ԫ5�x�`��������?��z-aA$ю+U�t}���	�gQ�&Tݢw�����V~@k�{Zr�L�������(��0��,�<��u�u"AB���][M�㝩}���X�Yx�KqK��~o��Z�T*��)�_�U0�) Ru�(��܅��Q�<��R�D�w��H��-���ܙ�.��r/�A�,����P_�%�'��&�F���i��Q�����(i
TL�>�2b��zP���"�P8���	2�p�.�� ���y�S��)��\a�56}�V���B�1�z���e�[��A�ԼX��d-�bμ�/QMF���(�w"g��p@���}�B�=_�e<�� �-����ˉ�ݬq����f�Ɍ&;k�+��j���)��'�^��vC`����x�Zӎ�Ҩ��֝L��"�Z������t��3�W���BGI[�I(����~N��=Cw���G\V�L�.�H'��(.��\��28d��j~?��I�N��<��e����r��nDY�
�Z��JN�>()��LH����f�L���i OxND6h��t ����w.%����=v�Mӕ��_���_�R>���u��9p�]����F
�OKB4�uye<�Q�u O(�1d��u3ŲN^$����_.��{M�s��X��v��_�5�O�$+�C��T�����h����hu���2�/æ�H��C8Xl	i�pT�N�Gı���C`Q��Ģ�q�Jc���Iiy����炋����H3�w.7S$0����)�,!=��97��霩�ʃ�Y61C�$��f l `��l�LH�dS`�������c��K��*�S�q��)�[ �ϋxvRz�y�7�\*MqH}©�o��� ��a'�A���|��*�Б�cQ+F��&�B��q���"�"�̓�4��er;�Qٖ�˧�4��cS�Օx�<���y��pNHT9�T-��5�n��\���Ͳ�G�u,a�0bu�rk���>7B���&N�Rh\	�L7PJ�#'E�`����̕j(M�����]�-��A��¡�Єu2�\f��$1�.����o�"�����5�>`��H7��(�!?x�\��z�^>�B=���8���J�:	}�m#����Yܘ"Zmjk/;q����1��~��A�عJ���b��������s_�ׂ@f�aD��hN�]������k0�J��$b���?_׉�i�7� ��qOW�`&q���p���%�S��/K|R�����=��F��H!%F��$�"Td����?� ��+�'!����!BFs�W1����d�*� B����.
�|N}��ñBׂ�y�z���|Z����0� ؒ��eT����V �'H+ڮׁ� ��}4�����Q���E`gA9���i�=�2b$lԋj�û�1T�{
����g(�;��L�ipgH��i�y��;�vdK�V���;�s6����s���h\K��/i����� a�D��:9,ft�ݣ{�¦߳�M���9�g,{U�k�v�֝����)���qZ��Ih����).8��?o�)Q�E���\��D�<1Z�'6���
\~�M��������BK`�:C�Ϋ�U��\A=�s���}��A���d�Ƌ$�7�6@6����J���b=�dYQ���|)k�*���h��"�ߚ�R�#�p�޵�\��3'%pR��4�5�P��(?mUvN���ҭcREA��גE��Q�)O�^Z����]��I#��2֬��x�`d�t�r��ιlĀȊ�o��+ Pkb�!��/�4��a[��c\h���"�~�&�7`G�#>���^%Z��gd�`���n-��C��샿%ԗ��(8zo�N�>���Œ[E�/$�@���P޵.�$�0��lj��%Ha�x����7�@��j8~�L�e�_ES�$���;����Q�N��-GU�H*��7()O���z�g-�G"UI���4G�.���˕K�w��F_OrpX/�d� (����7Ggz邏dc>̴�sq�M�����s�N�B�%2��
�C���[�eSx.P`�O�<W�&O]���� kj1o�
����l�V�0�:b[�.�=���Qu+��j r��Nw����L��8�����
{�7�aD9,���Cc?EZ�=a��K�'��ڞ�2�ϋ[\���%�q�#R��7�I�.=�����^��]TU�������;2�A:S�$�_�z}�G<	q�ue�}�E�$�/{JW̾��(�c���k]�i}�Q�-�)�%���' Ḩ��ί�K�3����(U�1|?R8"��b#6a�@i�ܤ�^n}��]��:,ep�p9�m��В1�>����U֮}�|�ǡ~�թc�6���X<O���ٜY�������M���c��X���I��}Ly�PP5��V�n(��.#��'\�ܮ�gU��lG��/��Gf>����#��4(�k!���S'�����PY�>��ʭq�)fڃ��c<oVB���3E�X�����+Ւ��.�|���40n�8`��ߦ�B���f����oB��\�pUj�EWž����׆�b'#��Ͳ�]?��/��p�no�PQ+DWX���M�����n0��l���U��F�6�/����-���C*���5���	L��ez�(BkK�g蠭��S����x��`���&g�k�u��,�}�D�>��TA��k���^ f�%_�z�QL�3���ԗ�g��qFԭ��~*����wi���E[ɫ�ʒ�Fh�t�@�~����ܪ��e���xM����V�('����+��y����zV�Y?��C*6��iM�Nm�^�Fa�M5b�#0�[�ۉ]�2���{�Ŗ��)-��}��h<&�?�U޵�Q����M�r?1r8|LF�7k�<���B����\!�s�M�G�����?%�Iko���Y~F��l�����S�L�
����e�5�0�!a�C�^HI�k�B�c�i�&5W;��g�[���GDMO��l�]�i;?���+ew������[ͯ��IhnRX�	E��1)�2~w���+�Җ�s�Q����rb7�:�ִt%}C��뺷;�m'TQ5[�ݽ�U��3}��/�^d�t'���O]�
�u����:%s�݂P�)�>48���-���ۢ��7e��*J��B�R�;� a��ցs�w�����e_�B^�)?�5�����4B�߂.��|��B���O�n��%Y�'�	��.^3�W�ژ��H]���6������rB�����s^���J"F%�5,d�.�W����}�M���d��;�`?��- q+v������c�b,�G�
m��Ư�Џ��]��eʯ���n �}N;�;]׼0W�@}ڰ�R���N閹�-9��V�� �����j�a�+�o�&'f�d���vjD�e�)���*���b�������-��Ҝ�gfg�9Wiy�ʟ�+3y�	����32�Ȫst�X[ ]q�Ы �\lh�������'�����'O�\��8e�.�y��N�t4��c��Ƒ�)X�B`m\}q\�������߁@(�k���NY3�^V�z~�̿�2_�jf�_W�J��O2'�����Un	�d|��q1l�ߡ/�r14n�8WbQ6?�4"��dD�)`��b�t�.eǔ]�-��h7y	�΀D5�k��-�����ګ��\C����gR�Ͽ���)6�3��.l�=y�V�T�O�Q��+dSn��L�������Q��
h��n'ǩ��/�1����br�T���P��<�1+�U/{���'�������+x@Ol���&���JN�(��P��O[�H4���v���"^Qt�3�͐;>I��V���n�b�`��`�^x�픧8��%m��P�1O�b,!�����lAl���J,w6���9�>ئ��-��SX���W�J�g�����&�"�����#(�AY��V�v�K7_�m[�H\��p(*� �:V}�O�4y<�^>��=D�Z��!9Pp��^_�����0ā�g��-�� ��V��yOjaUq�v���~Hm��������Z���7���8 �/��Q�Û�5�d�/�ȶ1������ �t%����om��]h���'L���~c����ޡe���V�r|$� 3GOm<�D�'d�Io�U�7���}}�%a�=�l�g�i�Y�R��&�q���T���o��ݜV��˪�Pb_'V{ǳ�N��Wu_"�����o�-N�&q������ٌ�r����0�[`�B	̺��ft��(��g��=�jy�	K��Q��LGi�ޤa��_Viz��������Z�vA��'gDxm�ܸ/�}\�A˧���\���)�$�Q�?%O���E�a�Ms����j�0�?���Z2%���d0��"�򘓱i~>~A9>�X���z�ZN�g�Ot��:�=6���Ss|�N_���d��S#{@AW����61L.Lּ7��� Ll�?�"?�]'����\�Y�:��$�AP��QH&�z:����w� N��zS���սe9(Q)�#씙0mk�EW%�EGFL�֚S}�c��p�Y���L�jQ\,��Ek��+�EH�Ʈ�����n4U�9.ZA�vuP"�T6��	�҄�y�	����ܙ��I�t��7,w����5A�ݞ��k���2(#�c�%�gAt����t��V/L�A�Ed����9�֗pO�{|2�g`_a�F*�ʨ���1ښ��b�ϴ���*�\��`�0��qM�c��D�f2<�SQ��\/`����s�71'F_h�]0�RA蕰�T,�k�E�鎩���#<��E�� �]�h�%���_��/��&!5R�?�5X�Yd��{����:��Ü�i�sd^LT�B����ND�v2,�A�6�a��Y[�i������vy���J���y����1_ѨbK�r?^&qy���~�*��ʲ �-.�����(�3��2��8t]'d�}o!y��&/��~?�_�����?|�?u�cG�m��_z���t�h�j��/X�ArIm��~t�E@�E�C�Y�e�D���B?m�;�
U��"��.qr�4H66<d,c����%ɓf��oan���&��s���ԙ}��l ��>O� &{n����a1��xt��v��>�'.ߊ��$��q�,���D�DUt�YE3���,!|w��8��2��ay�Fm�YK�H_���kg���j6'���˝���)0��c��A��MKe�F�[q팛�5�� ���r��A�ݮ�r���6�^V�6�`����X:5��dx��!͠Ƒ�Ɨ+$��|E�H�T���O>_��I�ɸV��A�蔂[Fr@���Բ*�~ Fycn٫�G��g~�T�P�n{DY�0�SC����)�<�Qo����pg�hpy�9���F����.�n�a/��_��y��ȑjzm4��B�M�4�d�T˲ܵ�&������z���ާ��C[�^�Y���Idq�����t�}�>��K�vP��s�gb����?���U>��d֌���.a��`5j�Ffw�.D�)g�8���u����d��_
�Y���c�$�|��:������"�i;�e�t2Pn	 �ӹkG #bm�v$�Yde@8��O��3���Vr���G�L��E(!���D(�V��]�4 �n���t��zIn�^���
^��@z����v[RZ�,�r`nd!��扨��ίH6��ΓP���	Q��ydj�r[��.��g�(���l��ڈ�\�<���ܸ���g�t�F
Գ�9�RռHo*�S��H_��v��Q�)���]0�\r���z��AqZӏm���<.";!G�x�	iɸ�&C;�>+d��>���X3�;�z���51�������P�ݜ��".�F@��R`��#���Ӫ �>`��.b�;$���c�;6��~~��jR"8/���RH�`	���0�1h����?4̭�X*E��W��6����
�	rǟ!�xp��('���@N*�\cc�S�~��zn��l����6H�;�vPR���=  �S������J>��hw��op����En�>���U/ ��WP	F�VR$LJN�f1��"�j'�Q��>��n�ڥ��Փ
�����;X�� fMx��ü�����;�9ۃYt_P����K-"�Hj�D���u�M��/L?V�P��N$rS͍�i揩��� �|_;rTlۓ�[A��1]��~IhX@q��1���jN������qT��L� �\��(}(�D"�Q53���R^jZHZF/KG w��Ͳ߀���u����� �������7�*�U����4��I;r���~O�lb��ّp�鲕E�-=-S���v�������<�\�(�uG��>,a@�7i���g����wl���������[�A�=��i`���$W(�G���^�$<6���gkKr��ԍM$�k�f�X��`U�3} ��$���z��2����O�{W"-�e����3�	0۝A�2�S���3��t��Y�2�6JP2�q�&�
A����������iv����MpI�[b�t���2��QÌ����<9p�N�;��eA�i�	���wo��@K�1^���K�7/�m8z�,�3��,3y�A���� �ϳ��]�%,�i@T$/����1�"��1_v+��L#�:HT$O�]'�:ҔpBC���MB�ӝv�47p5��.������i�,�˥���*��(��A>>׉e9ɕ!�c��iІTe��_�����U�3�Ϡ��Ò�Ì*�ן��6_�ַb�#�T�;�Ԣ���U��Ǎ�����sM���S	x�\�̩�.F��\3�,l�,�d
@�'�g�?��@ӈ���=�3�d��Z[/`CM�8UxМ_���ʺ('%�{h)[DNz�w=��Z�%.[,y9�b��dȨ�8&���O}���4�͂8+^�f���XLv�G�0n��P���T��#Y,��=fv2�׃��+.�1n@�6{��m� fg�K^�Y�U �*�T�fV��C���/C+uC�SpIډD�I�)IW.���qUk�7������FEΣ����ā��M��jE�tZY;�#�j����N�WEA����?�u͵��I�V���+�ɶh�á�C�A|�����zc�`AD!h0^����Ie㎍��1\M��!�_��d���h��Q�r���4"�`���gd�.v=�s��c�s�����}|a�J򷲪�F䂫s���j7��q��F/X0S8�C'N|^���bf�,���Pq;��
��7ԕ]>���oM{֧a���<|���v���XBn@ɿ��n�x���O^��HA�=S����T�7�2S�q�8M��v��CiCQ����6t�I-���,�C����$e������t�d�0��~�Բ�:<ȯﴒU@��U�92�5࢒���*F6E~���$�Q"u�:xӈJv*N�T<��7���+�~��
}��8���c�;��{i$[W��*�'�W�,]Ⱥ`_ɉlMk�B@��f�e5	�h"���� �r:L�d�$�d�ȹ�s�
x@/_���\�'�]!V�B왽�����+�u����^�* ��q;�¢Љ����z���{$Z�I�V��BC��C��nN��I�8��EU��*+6�AM��D�Qp�6Qe�e�乚�ƞ*9�P[k5}`4�v��gGd��as)ֈ��fyY�+	{	�8����^��}x�:��&�{ܼ�p�0�B��M�?9e�^�)N��I��uc�����*��A��f2�;?P�ơ�J�{ܖ0����;�E� |�^�&���9���(�o�H��7&�A��RKgl%���2���LNV���>����y��c�\�ϵ��HЖZ�����h�����@��������)߰��Ks㟒H,u��l'��ȓ� z��/���-e�
��3٧�|.�<W��1�߄ރ�r�1�>JQZ�{��|a�NM���ˇ���i���a��ub<T��)��r̩���h�@b�PQLo[��a�V�����b(dQN�V��G6�x���m�j��)%#\�8 fd?X�s�D��d`dg�Z�ͦ�WNXˎ[DP�7����v7�
`����t@�zc#���ZґB��UQ�N5�	�s�Ix<u�������	ꌹ���~������.���r�K�_B�]�{�sIE-v����yg�ï�iW6��v`�o�8�3��a����r����o��	�B���5�o���:-�Y���] ��m�ҩ=����
g_+���w;����Scmr$I|q��,���o{����u�@V}�禶`T��P�_a.4sʈ6D	�TI��0ۅa0-(����1���LBl�4��݆�1t�;4�j0�Ү�0n�Z�p�^���qQ�g�7-3x��(�,	��!/ ��m���gO�a�u��~Q�f{����u�\���g|�X*J�x{�L�b
Y�Z���1ʡUF~ٌ<y����c^0�4�*�Au�1P������!}ύJ���8��*K��;�+v�kcHf�3ˊ�x���9J�����RjQ� ��'է
0��rauU�QT�Sо%��������z}��L}��7���UA�������&��&��K$������	/�[��ewI��m;���8�:Y�Lχ?>"�>)\�����!1sY�v���Ay����G�CTC��+�%6E�����$������.�8�Nvw9ء��M��h�^Vu���gyCb��<�2�9��i�D�jKS�0��+^�K8�+�X �_��S�>ȃ�# �r�^���$aRn�ŝ���!�Q*�-�� r�y�tǳp��<x�a����W�,8���6��+ç�R
�(y��(V�
�Kj�55J�߱�f���z��4.do�uS����d�ʫ4D��+]�	�llL9�;��t�u�"FI�>����^T1�iI�+�n�%�ޔ�*�N�L�;��t鞶+��"@�5���L�=7aAS�9{�W����2ټ:��}/[��$�����=�+�#�1	��ZX'�ֽ��`�����B�]xý5�����a2�x�^���M��V�l�ll�M�>�M���E+����Q+q����ot�A�6 �����`�u/�XmwC%Q�L��������dO�%�	�L��s���6qb5�oi��z��0����dX8 E@��4��m�������͋�ǜx��������ybNL����¤Gr�w�s�E��Y� �7d���i�hz< <��3
��Y�D��3�ݽP��J�S/R���y��� JG��+�{u]`���NZ��lK�v�"�[kMW��NA+��6Ja[�	J��(F4?�?�R�#���?��qnE�[�M�����]w2X0L�w����hX�t�a�7��R�#G�N�DN�����v^3}p-[�w�d.r9�e�K&�.�	=/�X,J��p3� Z�]N�oI��{i��T�X&џ�UaQ�{�+�IK-�G��Ī�.}l��Y��Ks���,�\e�_�7��.�_-I����%*����<g��n�g"B|EMR��PVDg��T�Eϯbp���|k.lј��а��o��$59�� i}��z��߯d�Җ�����R&�����I�=W���g�}���O�7��"d	P1�|���]̺X�9Kt9�PB�*_#�4Z��� %;i��7�j�eU�����z#��G�9�G1�r�<�	����zĩ��vi3�+�S� q��X$GP��#��U��w���y�䙡hi�t<���I������J&�1��_�?��AC�9dŊ���{ٷ�C�Z�0�S�۬��"6�}����ZvQr�劬��ի�$f���o� ~3�����X�}ܘ����x��g~5 p��Nv����o�5�*&���alo7��j�"G��^y�?d�.�Y���?��+y��lU�lX ���LCd"G�P{�і����������%������=��P;I�&�QiN�R�{n�
6�wΠI��N�U��g����>T���Sh��	�t$;m�;�`�r���h�ϙy��o��D��I�\�����:�[����g��sa�EMJ���>"c7���驫�<bTc��F�PAB��ȇJI2��B�����8�8�~ŷX��u���e��ݎ2t�4#%���(�W�ᖟ^���Bཉ?@	��0r�A_Q�AV~`�Fd(w�.�(;íD
���ꛊn�1�d�}�oE�ɇ*��[���Y���?��\�_��'��KZ�o�㴪$�ѩ!��Eq����T_�2�X���9� eL� �y׷��d���J�� �������+�{�% ݐr?m����S����y0��.Q�0A��5�Q"(�3ȯ�3�&�˝R��k�� G���f-ԖL.�dy���G͏��I�_�
+5����`T��N�I�%��&W�e��ذ�'�͈i2<���a�ó)݌;�!\[?=�Aв���Ӟ��¸h�Ґ�t�ж���q�(t��$\�Ϗ���?�Л��]��\���?Vau��X�h�h�,��s�[ Ja�J���`�Y
o�Uhh��f@}I�|׬5`�2Sظ��0�Ծ�L��ެ��������n�MPjA��o�xZ\ܵ���c��|�b���)��dL�nSU?�j��%�+>Zj�ģ���ͳ� ��m�Pw�ٵYsխ5��(�"8�f���,����I��4`��o��]n���,.��QL�Mq��d�L�z����!` �)����X��?,�q�2b`'�m���Y�t�X|5K'1%E&<,*\}U��U�nm��g��M@0w�B���&��\f\�Rs���t-��fQ�o[d�?��=�����0��fo������"=���k/��6�E�7��(�qN��P��@�>���  �D��'E�B0al�Q�%�� hf:.���-�,�g=l�9�U{	)ϵ��xI�~���,�(	��,Vv���l|j�YJ��#m7S��!lC���X18������ߥ���[������P�N��D��7�e+���k-#qs9� 5�1tq����H��Hywm��i�]9��J��	T$*�Man��#��3��}���.���XQ���?GS��|جqQ�ZR�dX��0V��RE1�XX��{;쟽���m����K�ܺ���5�7����-��NJ���o���#�5�"9$�ì����+?[�i�� .��,��~ܓ�\�4{�[�@�:2o(��]�$�M�]O�9�����?��7>nM �x�TF�|�K/|E��+B�S.
��,�m.�I��~��}���r"�}f+t�!�RvdP���܃�$�A�6��H����s�.� �������82��?��7fl��� ��τ"���k�l��s�S��1��h��M+a�N��E�hAd�$��M@�089"#g���X	me͞2Q��r�K���i���	��+���6'�ݹ�yѹ��o|7~*x�������V`��~�E�0��5{�� �'Ȏ"�/�JL��q�^�J�w����R�INQ�
��Q��#$S,��t����0LYԹp�e_x��؜N��
Ɓ�Q�j�i�0ڠ������xh�`����;�sFXca��m�$aH�-�-�\���/A��£��R?�&N�(5��T5��R��2�|$�s�O�ެ1OZ/�[�; ��
��H����?.,��p�Z)\YL��X��!i�}�����H2�g�啥 {�2fG����Aܒ�X�5�c�@�ې>c��S�ppB�P^�1.(���"�
tmo�e.d���a�!~D'W����o`�����Z-�a ��={�b�eZۃ$���)E��$�x���`p��D��Q}HO-#l���!����.;���/�1A��@�w�yO�!��TM�}��vL�C��:�N��*^|�Q���7W5��כ��o@��ʪ��+��f�z§:S(�|��I��Q�Ji�*Ӈ/WZ�&8GI^����-�~�w{2W�O~�#[���Yc������j�5�ȡ��Su0�V��_u}���>e5x��	��=9�A\��0�ϊ9�^ۥ�~5~kk�\�Y�v���f_2�>�s�$�)�^())���?s���A�x�	k����"�/��q���x^jm�%�+}�FzI֦�}�_z)՚R������˯t��J!�y˿��J�"��D�'1����V���e!��`.��F4��EϼJ���!��{d�
�\��� �����������a^=�,膹����G���F,�/��`�ߚ2R��Xvo&W��"��2���C�r5�����F�TK�b+PSe�
@�b��j��p�t��lR0���=ji�i�N��ǡ�`G-�#��z �h�j_	��ס4��J�O��ES���J�W#܆J��̡h�nO$K|�^�����m�����R���H��^��YS�L1��@/0��Jr|� )���Mp���<s��[��=N����j-�����G)�s��W�ǉ��x��}��.�l�Z�E��m
}]~�.>D�Td��(*����$��+ҏB�rl�R��y(���DH@i�v��OB��s���g����}힄�;V�*3p�〳+%�<7�s�(`��rY��"����iU�[�gm�ҥ���8 �4ޖ��j�;Q��֨��g�T|�M��Rk��+/��h��@�.�ɉ7b�s5��n?G+� ڒ�sP�$Ѕ I�k5_�)7�	�Mc�8+-e��A/��]�mB1v����7��C����[��sG�о�*[1Կ�����#�Q} �1tk�ԡ9� ��	�V��_2k������q�������u��9�Q�Ҏ_\>�#�vd����=)V����;��.����7�RE�o׉U��&����#��O����2AA�]�a_w$	�mx܊��}�b����)��N��#oz�cn߰y�'e��pcВJ$V(޲�ŷ@�Q�^�t�fY��\RUu���H��q��2��ZF<9���::�>-�fYA�ͮ�Z�*���mI~3[{�n0�����m�!P_1�O�?4��s�������I~�e�9�x׳�u�3��ء'&����0������D�˷��~Lo��ʩ�+��^p��o�K;������t� �^Z��蝃DK!�3w�qCC$���*��&�.a�)/G�:���U��F���%VRu,��L�[��Ǖh�(����C�O=��1M��4�����qA��iԩvRx�S����v ��hoW��=�@��E���Ձ`�-!a%��n����x�\Xw�-.��Nt]
�0��M���� ���]q�H�o�W�d?���X
���uO:B���D�i�J.��\���õ�.�԰ud�b�@`���ϸ�JA^����5�V(��*��������0��ߌl�@+_?f�)=���J���JvEDN|^��g@��"C"9}W.
e�؛�%�]tO'�1�G�N%���u�R&��a��c̢��&B������&������Ћ9e,KZ�U� ��?��?*��]^�\�jZ	ͷ,�A|rH��?�0��0�A��lN�0=N��.�8��"�yi6�,V���ƀ�o�_)D(!9T��!3j��]G�g��P&��83r���p�)�|C/���De# ���Fެ񗉃(����tV�8D��a�_ ���+��:���F�t��>/+QZ�ܭX$����O<J�+��E���5gE ~��OClt;�(H�BMDB���&�RZߋ����?x�Hh���Gӿsg��$�=
bf�5�;l���%��E��7��*������bl9XH%d ��֋k�o}�j�c�Im)mQ:��Q��VQߕ�Shs@�E���wȆV�V�0�fp.���Ɇw���E�^��K9�3X��|����N���J ��D��[%��ط�_�w//���6~�` Y;�ի!g�x�q�,�4n��=��˩�v�'�;��Jd5(鱽x�⦯S� �N
�U�j�CE��@�����Q�N߳P�_�)��O�����4n{�� ��Jn���m�Ƥ~Q��Kw��#m�!e�bt�p���J�r˗PT���n�5@B��8�� J�ݾf�w0\���j��&�T^��*���*�U	��"��/�d$q�M��
~5u_5�d��C����>7T;��B�.�b,	by`��k�U1�^I-�g�ڳ�"�]�(M���L�oEϿ�d��B �	�; &Du|�~��w���=o2��<7�dQ ��W�r������mp6�� �
i��U0傎(xrMdd;R�Q���'��
T�I�H�[�!�nЩr��~�����jV�P�~C;�| }����2Cl|���=��C�  u)N� �G��ʠ� Rw̡�x�ꨕ��.�N�+¸g�j�4ㄋ��Ӹu�7�f�(�����w=�!k�Vi;�x�%VI�=�T��%�.��|$�&Q��D�`-�d9��	<��A��C��hE���0��*�6����y���jWw=S�g��3���5�k�G
O�]aG�)�7�6F`#kݥ�+S�@5$�0
�\ �NDh�aP����O��iZ����u�hE�������Ԯ� �/���H-��?���Lm0(l�����{�fա[A�����B �#׆���$1z����Z�H�:j��'2�X7�$k��_q�7�>Lk�@�% �}4t߈���̑Wu����j�=?��a���<��"�[����WZ^l<&�e��'�X��ch�FL:=z9��{F�LE���&z�_�f�s��<m������UD��uz�E���?��X���&"/B����2V��4�m������z���Z�9p<LF\���@�0]W��TY�x��5g��ES� �Yrd zϐ�%T���ik?n�3@��. ��W��?��^Z��v5g��!�%�31�+)��VU�Н��zV?��ŕ���\m>�4bo���з �6�w$��I�(����-RV�泏l������]�}�ƕm:T�P7Å���h/6!u'04Lܑ8�&,V�y���!Qr0��s�S/� �O���/�֙�T��@��#V�Q�s`Y������Q��.��?����,&��$�Ih�]�T�h�4h/��zخ\I����Ӭ-.9G��VgIt�nU��1�$oFۓ�~�-�/Bd)I�o��T��ҫ�{{L_l�_<�ʂ
��&���\���I��2vZ�m���#�(I���7��tl��'a+u˨F�6WO���%�Q��&�'���ӢE}"Y@��χ��_�.td�O	�y�;�Y�_)�t��7���~�G�݀g�ކ6���c�_�EH�+��ã��>�e5i����
8����s�88��D�me���W�ojה����.n��;
��GЋ�	���%��M�D�*B�Z��*1�)�����t�n�db�?��T�:A��{\z��fy{��#�|�yt�Fe�|�jBB�i��+�����	3�ԗ)I���'�rb�3V�ȧE�'����,�F'�b��G�~g�d��6ϭC3i(���pC	;���y8-�����٢"��t\�rO�5�Dj�B���E�0!�{�2�x����v[3
��IK?�G+P�� �˵Y Z��lIl6OLu�Mc|C\�N�p�}w�LÑy@X�nq�	?[Hu+�8�<���s";��S�s 9���:r����mz�ڮzt�;�+�����|�O��Uf�J�����[,h�`ؖ�B�R.�Ha�+r7T�h�v�-ITs"��*� MW۴v&Y�Q�n�Բ��&V�ļ}�sxwT�vI��6����%����l�\��]T�U>?��������;)݉ҟ�����g옼��[�%�b��6 8��v�&�x�$_���Tesi3|ZT`��XX[���E�(0��9�q�^]�:p�l��vB�p4�)'����iE�j�3w��7��a.k�Z5�����*��
(��=�g�\� �I	����/(x0�F�����f�q����=�'�E�,A�����z�����(,-��̴�����@�}��%�`���󘚆�@֎/`KH���YYt��oQ�Q��ɲ�u%�r5�8I�]���"�I�wH$N��ܸ��4�ׂ��������|+���������04ZzpQ|�ٳ�[s�v�EW�2���[ߊQ @��	ŎDү�+��.���Ӿ �[��we�z�Q4�b�
�E7��+�;�?�'�Д�c�ƒ�^=�E3▩Z�yH��
qJlW�ؼ����e�f4-��	�f����z�U>!������}z�����Zx�_m�K�P��x���Tʗ����ɱ�j�II�Ȩ*�E^��pp�����NU)��C�u��K�=�=����D~���@��,e��L�aIw@�kԫ���ه����|�`�@��<�r�ڪ��r1�T���6��':��O.�ܞ�9p
?�y��7k�3�W񐽻��V�p#��u������x������W�eo��S�n���|J�4���v���Vv�_��z.B|���%�b�/�l"���(�m��
�Ô��ī�@�b/�~����64 ��?f��PL�������r"�t��^C5&�ɬ�9��`�=`�K/x�Ը�t�(�S:�(����}�
}]̹7Ŭ�\��U���=�۞1^p���	�7�ֳ�n��qy�[I,�|�%�j��� ^���n��0 y�N�_���r>�I�֪�<�{$�j]F�s6�v-�߂PZF�����VE�D6�QR������ɯ�}G�E����2��P٪�\(��C���/2��k� $��&�M��P)3�����F�ۛq�qc�Mk�	匝�b����tm�(L'��[���;�?��R���j㏬��:e�;*.�Q�nw~ ݶR��J���]����m�'2�X�j��Z�H���l�O�J�R�;��2m�W�^+�q���|L�#��zx,5V����Xb��Biߢ�<��*�����b�g
�k���R�?#�w2�0���Ȭ�`�w�{��z���4z�r/�G����ɪ�T�Ր�弽�R�^Q�Q?m����+Y3�"~ɳu���h]��?"�t`��w��Rt�:��Pj��]�"�1�a�z�4�Э.��n�B��A����4����@GT`paA!�����_�4�耙W�1qgt��~Y���ob��Z��>�vi�]�K�0�RN�5ckc���&��Z�@i�	U����?(�җ+`�ѧ�o��
>R�[S��,!��Z�����[�v�
�K����Xyh�� T.���I~���x�f;�m�O���V.nDs��C�f3v&@k�)X{PbXDO�|�,8�i�#����)`]�v��.�&t�"_���������6.}�iyZ�������� &�t��=./�À�Mo�O�����HҖ��7�8v��>����H�
!o���G�����=v���xpo��n�U��>K�O�8A��י�v��tr���ōh�ah[��&��Q�̭�*Љ%gVI�
<�0A|�w�!�}z��B%I����L
�2�z�y��������V�K#�wP_��{�>�v�[ˑ��1a�>Ӏc__+"��������������xջ���"��9���e$M+�m�r�n0t�߁f����5^p.�7q�NCK�v7���m?�(��|��<U�S�2�*^-z+���7�Ǟ��/�r�ʍ_���--˸�Z��zQ��|����˨�ۻ�Q�ν��{	��>�5�ʬV��6��-S� N;��WH�-�q<�أ��P&l�s&>w�KB��fC��f���qY�лc�a�m�VaXóA�mF�H��L�\���	���ۈ�G�[����+�n���O�o�?Fk�Su,+(��I�k%b��X�Aϖ��イJ��S(ˮ�z}�.5B&sJ½���S�"�>�o�:F}QT�!���7)\�d��w�0�������>�:�/�ԏƧ�#��nSy��-yr��a�.k*���a[A�ל��j�"���j{;�[��=}�6��)�<�r�S���T��H5U;�Ͱ�p3���#a&��D��e�F v8�UB�{�;:���虌�=�G�u��x���}H��>���݀c��ׇ��8�F��7sg꾛c�)r�'��ڤH*��@�FOR�aO���G(�q&l=�n�v�A4�%�����ˏ����p:亏����jdݾ(?�j7M݁�k(�y�%~9Qb"��a$.���7SO�_���Bl	���A^?6GV`�Ɛ�<%#�]��2KkF�m����"�{� ؝��������N����J�{=�)� I�z��@~�����>���`��:�W�E�S�l�y��e�I5�>jz�"Q(F�~��ŁlO}�@�.�~�$�`�y�,�g���z�ܡמ�p�����=�bfC(���EI&�G�20J4��m��#�I��e����P�T]�w�a������N�R�i��!��P�;�"ȗ\m�"��ؚ�n���n3������� �� E"Er�K'h��r̅@�ʢ^L��0:ˣ`�p�iv��Y�)��+s@w2�!� �T�_����X�w�^���M��С��[�K��e��tb9�O4�'���Q=	���J�u���x�!D����t#���р��1B��	������Mi�Ü���L:JEg��`F��� �#5�[��v#"jW����~24!ۙ�p�M�K}u3���@O��Rv]��U?�J���Q$ ���3c�^�Ι������w�&��-wP�O�@ɔ�r���Φf��j�?==l�Z�0 �m%��H4V@�@��l�u�r��	�q���IF �LT��pw���"�n�x��m�J�g�ֶE33��r�θ�2��wLN�:��[��C׺B�������T�rJۻ����r�R�˅��28���2
�{������Uj9"�O���Y��ʙ�>��B	����H�q�:��\J�nQE ͺuj�C�2G:�5��I���������BS�3$�c�=?�����g[ YP�����c֚;�-@����J�c���p7N�l��e�k3����O�z\W*Ae����:��;#��?��E4M�u�C'�u�b��p?�`�O��M�Y�9���+S Z���`�~���/�e]8�i��{hsCg[��*�ȵ�\'(��t� �T���>[E���GUf�Y��Y�8���)tK~��1j`��y�9N��H͘RA=�B���8]�#h�L��J�h/^|(&a`�4(���<t��rԁDa��� 4]�1*����/d��@5,`q�}�O�`Oe1E��	�[b(B�x�r�O
�\2���|F������S=��W�_�t�f���R���m7��̷(d�A�v��K�底@=у�2{N�[���|�õ��Ķ����\H�Bg��&��s|S2{��ч��Dˈ8v���,�Ɏ�al���к)5��U�痓静��ѣ��k<U�H&
�I!����iF�5��4gI�;ΐx�%���Q$ݹH�|����_~[����t�1(�D��A���oʐK�I�x
��P���zۨ���a��tp@O�����Y%��l�2�&e�.�[�H�D�ozη�a�����h��#� ��a��Ę\��,��dv$P75�����;C��`S�!�$������R��֛O��bBƄ8>*n���XヽA��h�}{���L
���˦3BYp07�=Q�+�&M��m��V�VW9����y��΄���r7�pȞ�Q�?������~eWhb��'���-_��E�GtM,��D4(`I�*�SZE��}��4�۳t�1YQ]l���c8��
Ru��Ɩ�}oK��]��	�z�*QyBOx������`*#����A�S&uE�2��![C����d
0�w[�U_�?�-�S<�H������-�59�2q?�Ms2m� ��3�)o�|s�g�Q���,+/F��� ;����E���x�F��_5a�3����;~�r�8P�i�S|Yy5^�/Q2�7.�G�q���Fo����$o�Tl��lJ��?���?��O���N�U �l��gn��w�rF���HNt��r�X
A�S7��Twc�(���ƶ�qR�IO��}F�b�(�Y����3 z)�z�-h�>�U�W:��� /�)\�p�ZEO0}R�1���`�n���
Py���}�3�-�G��>���}�l���6�C?��Ͷ������L�V��9<pF�* ���c�|�}f
F�������a�h��X�����P<z�~����}�:�63�u=��6�w��HO� ��U�V���5�����S2z�A��[\�n�BsǍ.�S�ѽ|��eǦĂ3�+��Lz�ќkY�"����5�\�/�<0���߂�1��������Jg�*s����i��N�N�D�0�<� ��ee��ϟ��1"���W��Ȝ����Lm��#��Kҳgy���:���\fE���Ӧ ^����I4'岊L�9�*�����+E�_h�J�R���3���q��fr���XYB�ԔL��z�7zQM_]�	���2��ؐ)Bg�O��`<�"�H�sveu��*��G4䠈��$�_�
l8#) }�����z�>��SOǀ�^��ZC����SbҜXSaGyګ��7g�,�Xݷ<���̴J!��d�Nl�g�W�k8Ӂ��r] =fw��Y�.>]Õ����tn���0V5�@��@��i�P4ٟ��W+�n��<����1��+��gL��,Z���1>���@���~���I�$�l��	!��:e��,k�ΘtD�����������&��c�6��֡�ÏEi���؝[a�݆0�䞟=��I�۩o�u��e|���KC�/}�g���=�f 'FQՀ�?�oI�WC�;����M+��Q��'��'�P���o^"3�&2�JS�c/ni b��<�2���֯<�eݗ5����������8�j�(h?��,��d�4ao��Sn8�H�aF�V�W�km�2�te�'��F
���:���!e��v�_[����bE!C������H�/�4�-v�f�ϡ��)�1�����+�����.��WU��u�sNv��Ռn�.L���c�MȂ�y-�By�c�����[�cʂ�����7�mB��|�LQ��(�V��M�9�pI`Գ�L��c�n���H	�'�y�/G>�6Г)�ǂ��zm�����3us�&���ls��ɕ4^!RS�@8��$.jT������Q�&�S{���[�����m�@��׼�/F�,�c�4ؚ����@�:U�)$���E���C���$����;��'`J��`J�	�?=�� �!u2�e.�?�&ħ�tF0b�t��<]@�@�2���嬉ku�'.�N����h0[gA�� ��aC��3�j
�-�|� ��u�4����pKhP��q&O�9S�*}��F��6�ָ��X��$�`дw�f��w�$�N�din��rY����Ժ��I��Ã𢽋�<�����76)��� ����,Zr(Wy$b{��冲Y�b(C�Ť���(C2�(�eԱ %%�dW��������?�~��r��:ʩ���*�z���%`c'����*�|)���V~ƭ6��Θ�-׻x�	�R(o��uYs�����,*��+9w#���䢄������ɱjcΰg*4	�w�{��h�'g+wAT����<8}+~<Ϥ��'=�Z�4�9��?���p�b�R��΂�P�l�.�41\�_����Z-��6��5���t���+���lɍ�̒2�! ��0�۞���`�>�^�-,�Z0�^��]C�7M��w_���z�( Jo�+NN4I�!�9#�na��H~���BC�R��hU�Na$�F�I�@H&�讼 �'#�[�4!����v�!�~�� /=���J�I/�i�U70�4Ԙ0�Hk��:BL��V�����N%@��UǊroտ��
��<#���_f����)�O��S��[^83x��L�18��9.���ϫS�K�'5�A�Ɓ��:[�!�`��%D (Bߩ)j��m��oq4��_I�۵�1�ho���OQ[������x���7���*�v���y!%�'�z��Ⱦl����Ī�D |y��C�P��eN\�c�E��|��0[i�l�ֈ�ޢ�L*�*H���׌шAu�S�����[o���&漊^K�Zߡ�cp���WI�G��)�h���YG�`�\,������5㉳�1i�\�X
�����75��l��3V sYp|��Y��>p��KA����$O@�AQ�Q��H�[h�y��F�jh$�J����:[m	?�!V+�Q˃����[��I��6��h�}rx�M`�ᓸ��da���5wO�J#��=RDo�k��`��3?�d�ҝ���3�P�+��uS6 h�.�f���TK��y��f?�.���� 5���$�H���?�>�<#���p=��A]����'*˯ų�������MDν�U�;E��?�	�d8�尬qYs>�
Z ��bH}0NT��my),Ձ���Q^"U^�j��u 8O����k��x��mzFII	C���u����|k�
m	�(�ĝ�VR�R-���oXR}\���א�U�z2�N:}G����ݬa��=DSot��Q�:5�U 5ވ��jۯ�������[4s6K��r9k�"�n��Y���X�S��G+�>����P��������=�JE�f1�!��y�f���IR���zi�{&L����nՅ�D|���۪���m��M9]J�����Hl;K���1_݊�1*��減\;�J��~�IV<f���XBm'������+}�Pi��[?�����|���߼��1.L�xT7���JLT�!��V���i,�P���B%�E��8i����,�3v6�s�4��7� ��ò��Xt���%�΢=�8+2�}q����L��e�$���	2�@
�F��ݟ.y�-n1�o`:�c|s�gu'G���+�}J��B��j�H�p�(2^v+{:V�~�~2��f$����c4z�pr��>"�:�bo��݇���w^3𐪔�|}�z9��ӭ6��*h��g�%Աf\��~���˗���嫻��K�cu�4H�o�25SY���:o_�s+^S���h��C�yJ����Y%�N�5�x��o��ke-���AK)��`��	V��hv��>S{�F������6R~�k���N!u�~l��:
�����~�0�ιE׍��^�, �@��u^��$�~}
�w����s-�c��5z�h�rh�P�xa��N�k��K���Y�Gn_�c^�bbed^�^w��y�%���b�c�z�0p�E��E�/����l�K�|p�_?EX-�0�Q�s���*��$��g���m&�Nrɱ+U0���48��f#���2 �^f0��`�+Z�])��o�w[��}��Vt`H�8êq�Xh��@��ͱ8���dܕ�b�v�LR��%�&-FHŕ��ht~��\k$)�1�[z�"������C�����^?�
�;�/t�~�"�[΢;����s(9ս!@��	�ܟ�x ~�b��k�����h�����u��!Y$蛈�&_Us�H>�Q�c����Qsَ�Îy��H�H�s��T�{���A5*>�r��K繌�+�(�!�d������K�O��ڵ��mHHA�хq����}���&���LjM��1�j5�12�	�5e�6���@�3�I�Sq0���ȁAB+҃1�88�E.g�r�b����'�%�h؄"nt���bw�٣�U���dP.�����#�l���ؘ�C��������<�=��e�L�ծ�ą���Tp���8wY�rW���ޟ�����{����OM`��]�l���}M�������!��I0#ي���z�2���$Òs�%vw�������U0NQ4Xɉ���y&kߦ��A7=�U�76��f�yQ7GO/O�U��Dr4�(���(�N���o��9\�$ł��u��%4�dQ��F���QL�g���Q�(I�θ�j�!��v\�&k������:�X�ʐ&�[e�G�֍�0� ��^o�L.L�jh$�%�W����R��	O���ȣ)Q�>�\.?i:w�JyJ����%{�p�yh���`�8����v���C�u����>¼e	>���͒����%^�s92Wm��i���>b_�+J�P3���D����r匉��C��c�]}QQ0 �NΠ�>��<y	ڵ��x`4�GT���;f:�mL/2��B�z$���m�b�c��H,�!c�|�7�o�5�U�e�`��r�'��ۭH���=h�i%\Jc�þ==!��S=�=J\bX&�/����rUX�L�&���������U�q�_ã�����ސ(�[,cJ챕ɈM�&$��y��I\���^Z�dơ�j����g�-14�݉~i_~�vpk�A���; �rཅ)��ME�X&>���yg]�3ܬ�bo�Yv�;6�@�)X�PG�ڢ ��`͋�߿�%���~^�c咧�n��bD���}�ÿ����r-O}U�F�'=x:(UH��3�;|%�R�h�ٓ���9��	0iݿ+�	g��+`���5��k���R-�W�U��PE��f��U��ӣJ�jm�쾸��4�h�Á�̵�K��r�k����ߨA�u�}���C�UE�%(��&Z�6ˤ6�.��*V^7�ށ�,��L;��p�ʥ��L](r����gs[����m&�V�d7N�K�Du�9~T�����rs�B��Z����y� �����>��a��'��kE��l#B\��c�I����`�ҠC��_J���ˌS:#��uc��Z����fb��rg}?#�J�cm��vx�A.��C�����z�������U'}�H��#<�}�:��;y��$e�=�3���X�wMH��8�<���4[��������qL���j�:�j$*�}��Wm��wZ"|��".å�e�uR���C��񏼳�� :�AfJ��K/����ǥ�F��j�gt�7�
�2�ӈ�Kʿ� ��lě�pd��Y@��x�s�qW��*�>�`1�*#ܤ|��lۼ�n)OE�?aS���ov
J�!�`:[c�K�$*��O�����ҿ÷�r�v��	Tm�*_��|/>�n4u]���	��))�wL���  A��]�3��N������9'FE��H<�nGD�`�3#���.t�4 ��H@�A�Np��4ۛ�u���ͨ�E_Dl���x�,�p�;��je�Â�v��=4x.��yM%ƃ����;�&�u���ms�q��z�R&�ۯ%�R>�~o٠&ef� ���x�����g��7�����p+@i{��*�K�h	������G��Rq!�M��L�9�0�z�4>t(4N���L�\��Urm�
��c��L~�ͱz�ލ�+��x(&܅5p�r���;�~����ф���K�%�,g2�hnb۹��$�1%�A��,�D�FH&	f�H�-�X\ƚ:�)[g_�r��S~�Δ�3Z`Y�L6��}�Hc�"N�ʶ�rr��� �`�����@Kf�@����Ka�W��'4E��Zf�6	��������X�� 0��p�]w�2�D_�*�Ӗ��t*�Qnq��ۧ�4�X��W���PJ���m��E�*$��,�J�ľ��J�r���ĉ�~n�5�뱤��i��t�y�R"o��0�����,B��1��ԑ��	���N�Z#F,Ǐ�/p�m\�f���+���k��ݿ�_��.e S �N����Z4�����*�Gq^���}�R6f�H����h��ԍ����wq�|�w���w����m��8C�x����*V�p"�[L�����c\a��.�Nsp�j���Z����e�O�M+���z�=��� ��^#�3�l��9�4��P�㓄�������¹@#�1�5�˽�pP���JRp:�-C'�8��ux#��R\	Ҍ�hk�q@�'�w��5 db��G���l�9����_ �� pzF�d��TΣ�,���¶i�1�0�6��a�a�ߖ��jpr1k�8�R�<U$=n�Q�+��y�#z�ҧ��Rg�����!�!C5h�|G�(�`���)���\Y�,/+�q\���t�u���'g�Z�Q4��M~G�gkk�.�"Nx�F�5o�o��.Л����n��i��� CFi4�]��S�R����D_���~r�P�`8�s����oH��&}���ʪ��u�[=�9�aڀ�O��+�C{i�GX�F�4���UO��� ��>����z�Cs88�'w���f�8�pےσ����N�I���R�M9w��x>cf~2?����E��8ek��^��첮+Vؿ�����E��-���E�4�X����<s���P�v#,��c��d�LGr�MH��x[���x�7�G�fx�q? |�SɵwEb<4�?��������nw�>^��׹��I-Q�[��O���E�dJi*���C�Q�)���|��iǁ�l���$=a�K9_���:>�f�m���s*	��F\��������T�⼣�eK!�S������,Fo���s���!=m���/N��������{#�4��W�g��L:D�J'�9�J�D�V�Fb[޿f
�wqsS��:�v�sQ�H[�9��\<nf�냨E��HS�w�))*��� �]���_!�_ᕱoE[?�H�CuX�BIJ��< IYO���|���?��L��n��Jb9�czU1C�py��͆8��|S�} ���}��2Nڂ�( k#n�!ZP�M��h�.�i�8NM:o�9SbO�	��.�v�.}9H�_ypۃ5����F������%���6�Rѳ�`�]a�a�zCZt�4�b��_�����䣙�Q*8�z�^+2�rU���������	cK��I�^|�b�r�o_�FT�n���:�!�nF���G9y��ռ2��-�FF�2B�����mD"��*��fG4v�����նW'�E��ӵ��SgoP���>':"���ܣx����Y�W ܱ�\p��e��J�s�:��S;C�[��ܱ�{l���~o���1��9E�M�|L�r1�O���Xt�u2���\����JHq��L��d��@
}��{�߽����/]�._(^�j�?��L}҅p���o�^`~
����v�ʮ����ph���L���"� ���A.g�V#�m/nv�6:ں��5,p����O=��=dP�ޑ���]�@�����aa��d�:)n)+�S�)���=��+�/8��F���wR�&����Y*����k.�r�
���OP�Ja[��,bls3���k�ܲ��Yp��)�Vcg�`�b&~�޺�h�v��HuS��6%`���8�@�G��3=�k�1���x��#}g<�x���B`������:��|B�Y��:[�\��,�����4����!-}�5��
�#��;i�j��ό�.�j��E�,�� ��_T[��YfP�j���;�T�y��u�s�3�9d��%l@���Q�XS�j(�a��'O��#��ѷr���k�������x�*�cl�(�=	m��S
|2����2���z].2����H�yt=\n�\�1�����Tڑ�PZ(*�`�i�D�m�TV����г��zM�1�	��޶�
��i�r*��q����S�v�d�E~�J~ݦ/<�wz�\�<��&M����$�c����?e�)��uS���. �>�(&�/��%��Q���#O�C3΅j�,����k��}�_l7�2+��^��kC��i��)���,~2*^�R�i�m\��jd&ogجú����ύ����K��9�Pc�0Ql��U��벍�������wo�1�+��#��:�+~�����@F^I��L�6
��]� ^���s�@��Ϲu�3v?��ĕ  ��5=���ӹ����bB�uL���^���>�x�:*��VgyO�-�V�:{z[F�e8��	�2����*�	���'O��^[7+R"��"Db-Za,�O���[����I�s;�p�g�sv����:G��\$U�����	�م�d5-A^���ݳ�ð�@�䕑�X���ԧW.x'[5��t�C�M�����G��G`2���#S~�9���1M�������L�����t��wk4���u�ajPU��Z"%<��A���8L�(�%i�%�Y�A�d&�&��� ����F�������8	��H)p��̋/�Ơ����y����#N6S�A&�R����|]�z��!RC��������kٿ�͹�S�D�7��r͛CY^�r
R�9���H+g�/>��j}��{���2i���Dҍ|=�ݙ^�L�j/ =V��f��(�&@��b���5t�X���ޘ�[̓��L{��p� �U���u!���a&a�d�ހ1���RL�V/#V{�<���`o�ě)ȵsO�-�(S�����9P�KZ���r�����\#|,P�᠞���Âf�/� ���g�M9�M.m�'����S��+|�Փ���a`���f�/+c#�`x���JY���1��G�aծ�*9���aV���Y 5���zRQ�'{^CPx�!��C��7�xT.�1x��x&Z�w$�:Gx���݉; g/�D��%g�Փ��&����
-X�꜃w
�AL_�	��E���`�2��F�<�`��ҿ���Nsy��ުx+�A*-|>�Ҁ���ga'�ݵb����O�	o����u���A��Æz�K��GKؗӧ��WW���OW�p�1tdP�D��+zW�T0M�d3c�D� g{/�
DH̢�!�6m���m�w?_=�Q|9,gaO}���i�$sN2x)W6�i>���m(O�T�m�K[�U�w���]gi���Ns�Cˢ�$�u-�n|/gt���L*W�C��Xh�3�bp}j��ѧꛢB�_"�3��t:�kG�������Iz����H >��|�_�ɑNf3��� �o��;��ӏ����	��Р��S���C2����T9Zs3�8L�~�]&�N��&��~ԒU>��C6W���vk^vFd>P!�VC�ކ�ғvِMoN
֛ƜrJ/+좱77���Υ��'�Yf:�0���>��؇��q�/�����M��U�9h��#v�E� ,�8����c7�XA�&�k���^����������A�6h+j�,&)�6��4W_S���E~��%.�_3��R�BgeҢa��9��U�BƠ�#K��A#�֤�ih[[f>3��q�vM�;
�Jͱ����v-�hS�=�?�[:������[i!�|+ā�؊uu���w��zIq�k�7_D���g�d3���Q 0/ˍ[?��t+��;8s�y�	y1m���PL�eQ2m����*�jADtD���;�Z�����I�z$	��P����\?H���Nk͞��:��2�+��x���ߺo^��i�ѶǦ.;j�A��(<o>�1���V�K��p�h7;���w�
`��jA�9�\�� �Q�}�%�W�b�i0��r�۸h�*��:N�&g�D�iq�ыZ6���8G~3�q�6$r,��o�`n2�2���9��3�eA;��ȶ�i5�H
$����Z���B��l���*�乄���(�<���	�G�$�$��|f.���*O��tFmI;� �����G5�	I�O+���]�h[���B����R6*���6η9� {dFRQ���e�FS����Ӊ8(�;
����¦�2����"�`Qez���6&�#��%�ٹG����Mp�GH���m��L���z���`j��WP�T�`�t#Մ_ڂ7����AL�`�*�3K{�P2�W�`���j啾a��*MS��� 7�
����5�"�(�|m���`��T?S���p1q`�i�?qksy����D��K��;�G�������8n}�����?�ۜ@	(�\p��R�~ol�!�U_��,��J�K#X�<vI��n��7��V���1D���x�>�7�פG�ɞL���	�UD@糾'%Q���GF�X�����A��Q��h\�z���ض��)���u�^���S���5�)d3��/����,H�G�xWF/�b(���ۼ��&���u�8��q����h2��n~i$lS�yEH�G�C�Ծ��?�����%�U�՗܂�C&�Zz��l�!y���:eߨ�&p�3ܞ�X���G*))@#��8�k)�ӸBO�	��p�����?ݒ�+�@k�Vo�k�5��wm1�-I$�����>�Kt>�����!T�b���P7� h>i.@V�~��}�f�1��)17���^�N}��3�'T���	�z�[�F�ޯ����g����56t�1�G:;)�l�{�����9���J���㧉��(d��`QKQ�7���N�ҽ>�U3�^c�֣z����$2^}��z���Ȅ]Oe�R�k+���+d�;���LH�g����zU9W#����<w7`�!�ܴe��8� �&U��9j�J��Ѝ]�V�^N<���]N�3���lh�a�Bx[]F]�k�D1גn_&0�փ�߳�?,�B�g2��H�k��M\e���m�'���(���w�[DB�i��2�7Xr�;�mg��NB�� �\�OI���>ѕL
�zS+(��J]o�9W��PR�_�G�iI���)�����=�J���E�-���36�UA�л>�01���߲��WJ~�%�F�e���z��`H}�L�c����w%Ic�;xW]�������-pS�����0g�u��0Ǥ����9:1Y3��_�I��8�\.f���Bć/?�qB�gw��v��ݿ���ۄ��ۆ4�36E�#5�B����L��N(X���2�f���;��C��}�[���F
U���pl�4Q��øg�~���]HP�r��Y1'�ٕ`��*ܱ�;�V����t���	Εf��8��$NpgZ��Z�m뽇֩���[U7f��=T:��E�	P0���|�{8�ۣyz��uj^��#>��޽y�U����\�{�}G�c�[Z��;��
Im��i�������~����Qcw�����p�7\g.�K��3����X���N�n��ː���f�s��׽��[��ĝg�.��Ax�?U�`wۼFh�t�`s7=x}'卌s�N��O��N�{iWQ{a��A�M0���\ꪹA:Ls�~Q�
�'�,p{;`��{֛	��ED���/L)��1?�������P{r��N�ZeR4�;:����<Z^��P��(URe�>&��U����� �Y~���l�V����7�h���0WnRb*�­���Ўk��n�Ʀ4�PI� x ���Y~�"�Ab��;Z��+%라���ͻ��<�^�M�6@��]�z)'��
���º�9���:ʔ� �/ ���;�o�h�ԭ��¦a��{��`�}BM
�BCI��4��"�q�e]�]�+����<���ia����Uv���{e�Ԟ��5f�Ҳ9\����HAӻɪ\y}�t��U��'�i&f�E~�����lOl&	���! nb}����������Բ��� �j)����\l�z���e���?}P���+�y��,1v~g��Z؈��c ����_�z�Ai��k%:]ǎ�s���Ă���j<�Eɠ
Ya?����{��]B"���B�UaȹJ54*h�� j��f�U_l:��x�qgI�Fn�Ȼ���������{������l|�M� ��N(lo�_	�*��2}�q`�bO���|��3`F�U�pn�K[����$m��j ��}B��"B��Я���₰��_�|�)OrD��}��Z큧�(-Bz:�LG*��5����n}��+n&?����e�?X��]�n;�3 A�|>���%�%�QжXdB�l"憂��(��" ~>�����Zs�#C�q�9`y�ʆ�������"���c�h�ﮖ}�44AL���b~�9�b	�.=έ���hS3\s"��<��B%8`��L�Ī��yd6��DZ�U�c �+Sre�h��:��[�>��[$>����]��M�y���@þ��5ʜ!
���ٱ*D���1=�X���B��9Z�BgG2�do�f���Kf�ū����z��5Ը쀞�[]�s$45=W��s/��Ԥ*d|�7�z�\ q `bEJ/�}���ַ�t���(�?Jp[����d'�#�F��?aѬ(��;z@;��(�lפ����X�����kJ&@'��Em��\؛r�c��P({Nx�6>����u�v�������Q�Ҥ�5fM4�a₍��a=Dh�Li�����K�z����s܎�Y�2�a�O���j�hx�Ǔ&�L��ڱ�<z����z�3��ǖ+b�� �03��_����]\���4�D���\c����,S �� E%t�Ѩ%ȿr+��r!ʰ֚�Wh��_�Ǵ�d��ONl�� E�#�L
F>B�K5�fD6p:���kV�u��?��K���K�h���v�"�͹��o�C'ӧQ����o��0~m�+!��� ��G��]�;m�'�3epd�A\r�����T"���^����L9V?hö����q�4�O�T�c��|���%��hhMp��/P4H��Y��4xz���؛G�y�+dD*\V��p̴8�j�,F�I=Vp��Y�	3靠��(�ݴ������-���̇��l���7�>� ����eg,���H+�c�y�Ӿ�7��mG�����.���(l�m��S������)�T\���
�l�Ѫ6?����a�(��m��R. G�m��e�<"�Cy�\3�߮��ˠ��qgyQʔ���X�����s�d�e/D�#Q�����7P�Z��l�Ψ�v�O�t��eR��l12WaT�|3��|��_�P~{S���_/��)<���X�Օ��.����W��-Sy�KC$B�<�ڌ�$!#~��G<��u�J��'�Z�H2�T�ӳ§V���f���U�{�Dl�^���y��@ˍ�\��kTu��}lԢƇ'�M����m[��@�᠎��F�zm<f����wM&�y�(��N`V��7�����8��_z.\cLU�1O}b��B�o	yEF���k�c�:YWQzGI�����7Om�K0�DS�!�z}Ls��@uE\���2���-�O���!�}wl���KB�m,�E�Ӻ��e)wO����Fj��f�P�;8@��<�3��=V�m��M���6��Zy~�-��ǀ苏��i�scn��kpCJ���8��"�r� c3��v��V�[�����nZ�!m6T������eA�ũ�Z�C:���@����0OڕPo-��|�ZY��ć�/�����NWg�����U,�G�:"�U��y�nC����؁S��m��
jFk;O����"�����q�"v��Ð勵�B��ٱ÷�/�	�++�:|2�(#!AavT��=e��b�!xc���;�[�-��>�w�x�(����f�~��|O ��Vɇ\�+�f�����C��H��˂��}Ԭ?�cfs���'���D��ߓ9q�,p�𜠾�%��E}����doh���
�:����n �.�N1|�z�6r�7Ɋ�fI��Zg��$?{����6��_��I��f����~n��H-p���a�-ä�E\?F|�sB�f� �����M${sx�޹��.���(�����?B�4eb'=F��Srg3Q&��e|��z"p�g� �p,��f�):��H�.g$z�/2��o�='��;l����� V�Օ�Q�r,��h�����N�'b�{���
���<���X� ����4,)|A�@>fšn�X�H_~���!b8/ӽ��+�RS6h�t�F�4�/r��C����6�sZ���^Q�1&DGHcU!��V��Q�*^�a����i��s1�+E�jΥ�r ]��� �,�Jr�V���|�#0R鎘��A�������@��=�9`, *p�Χ�B�����YA���!�H5J�T�D�T�,���{�:��ae~1�L�*obZ���l�ف�~�u�E���p�5Z��%��Gq8����ی�.�
�B}���M���
'��wo)@��j	�"�M�Ko���2#�+HFw���8�xHt����)*��!�;�b�O@g��7 D�=���Г�.��H:Ar/�כ=u
���l���D��n�ў�0�mĻXp����#��JEC�S�&�6&8�|�YŘ��碅��Q�syը��N��_߉�����x����؉�F�ý�&��V�����XR`��Noˈ#Z�P��k�8R�m�.t0�I��݇�P�Zh�(�Uy�9+���]ׄ5��Ƨ.'$�ݤ�>+��MƊ��L�Ѝ0/ҝ&�DI3*d�؛�J<��g�HRv�Z�2������!,�C��ʩ�q������n��Ub=�*D
T'��Y#�j㔭�����t�[��>?�(�܋�8�(��[5w��_{3�@��֖�y�-����b�z��3�V��Ԥ�����5QY���(��[�,�P��h��;½{�1x���	f�}Ryg�(��2��g��&xm8�	��ɇ#�6�������%��[��.�ө�v�j�

܆���0�0��,cY�9:����Yk����78ճ���2ń:�
<��.�")c�	�a�U�Y�a?��ж.�^}��-bWo�Nq�E-�u��>�X�}Vl/Gw@�����J��` �hXT��j:��#�T͚Q~�=���Pen~��1˭�B�{�&��� �D	ǽ�n7�2��<��"�;ĩڟDy)7}�.�*m!B�P�=�&G��R��y-H�pa�mo � K�u�� K���E}�>�@�&�;D���"�(Y�)e��htf\� {�D>���Y"�h�s�it�Q���4>�E֩��&��dǊۖ�[w�&d6u�+�Z�_E(��'/�~�M�u�<	�q|AR̄�,�D*l�@�o�A�A�%Y�b|��O�~T*Ė��������\�N�H��HE$���ɯ+?o�QI��8�/�IfhN\QAȭ?>k F�PI�#�1կZ����wc��  ��*���[7Ejd��"R��b�6cQ*����Y�x~�S��5�b�)��)}Z�,I'E#�ҽ?0�M���[;�7
75�<i�Y{�LSV$�a�6�ų�.������5���|s�(`�G�Hl1b�KpP�_G1�]N�o�c"(
W̐B�3�=���Z��^�p�!��q&�+#��Bds�0��v���0u혽v'0�ISz5_i��зM2�c#�%=�:��8e!�˧lqse�3w[���ܧ��/�swIc�r���i���(��&$����Y�U��<$�U��㈺�`&:K�����
�f�e^��ʚWkY�C6��8���Q���(����KY�-¦��ٚ��`BNNR��O�QK�U>i����A���
��lE3�#�m}ԒG�A��l,��X7��}��]+� $���uB���wΥ�s�߇q�ejs�n�BY.�J�vB�[��l:�g�"5̎�EM�w	���J�4h63���Y	�t�͗��z�c�w�0�C�Rn?/�"�0�l�aj�Јx=��fh����@��lZ$��#��1�	~���s��8�����\�H�|/���o4�,7�I��b=���l�L�e1���f^�u���ӨDj�L�yg��ȍGH���.t<Fx;���	:Y��'�zOIuN��]�^82��V��|I)�u��g�l��1��6Y��������l�s���x���:�˘'t
�[n
iW��Y-�F]��C�"zz�Y��E�wm�ȫY)����:��E�UU�I&�O;���M�GE��x� j��z�{�֟b%v�v,
��Ə3/�F��qW�������_��&�y��O���ώ$�<�_���[p[�H�d�>dG��5i�#��$��+�<�˜~N������xC�BC�sǧ�V ����h�p�:�Hi;
��Tv"[��ׇ'��Erχa�4�����3Ӄ�x�2�<Jv���"���"�	��Ӗ��z9�������	 F`��H��M.A�,<K�Fp���L��'/��.�f�[���k1ɦ�8*Ebൃ��}�m)0S���E��H%&0�9�G]Cw\��~�n���-	x�:4Ѯ�@�u9����i��m�W�oS��H�s,!�8
����A��ݣ���㵆7���ȷ�����jv�;La��,�/I���m�p��T.�$��(��BR�� J\ ��������Cf(��N�X��Xd��p�9���Wz���|�"Y*<�IHg����,yaFC�i�a�`�/R�sZ�F�- \{��qEo������xI�����ҕA�N�e�*���z�"�}m�N�?��v� 5��?�`����gj���3����ܱ}�X˸�8��x�q�vՅ��L�sj3X��HD�c�t]��J�l��P�'��N[�3Bdr��|8�f���=��l������Sx%e<��T�w�Q��G�j�nt�<��������Q�gś�·o�~F�ό���!m״ti-��a�Aחy�ļ�GZAv���icѣ�mҐ����y�B�O�C?a���o>�����$q�,y���4;�G*�L�����b/��h�݂'�{G���i��91ǯ�y��Z����K[�����l�w7+γ�9���S�΃.^7v��ޞ��ߺG�c[��`XA�5��x�h�2a<UF�n��~ń�b5��Q��o_x��?AvB����lh�U7��qnHD��G�W҃{G_�'�A���C�z"�C�{ ��Ȍ�������5b^�g:R�"�G&�g�1��s�[��.���2����]F��/;�0��-��y���Q�z֡�	w���֟_����0��Bor�F�7{�f9e��ֺcGj>�"i)�9�)���Y���?�s���\��ǝD6#��&��k��D_IwG�v	���@:�o!�71_���D>k�V* �~��UB3�|j)��U4�	A$��9�JGʜ���u�J��>��]��@�	�럩=iJ�v��b�ml��	���NxЗ�a��7�f����`=��t�n�$�T�x��u����;#���-|�G.���a��tI�����8����{���B�uaPZ���e��W��u=߮cj
�����pK�<���h 1ryx �]8���"E�cpD(k<=���'��ZQ��O��.N�y�����Y���>�\:T�ʝaT4.��װы[����/;�V6Iʬ�b� �r���У����~���c��#a�.���y�a��;)$����0^�ײ�Oo�ņ�E"��>�yS�Ґ$����Qe��f�gJ>����p�h^�|F���� �d��V����V3�dc�9,�`5?�]��.�,��\Y/^-Cƪ���&��W�g���<���l��j����hƗ3Y3IE,��OSzk�� �����Y��^�e.�ʁ��qҝ��	\�U����ο2��^�jA��UPN�*v�\�R�ܔ���Z*��#Ѧ/3���%��6l_�~�Kh�k$(PՃ,y3��k&�C���fw�k�`��}O�u���npD�4+�J^*�CIVt��Ә��w�K��+�� ��R�M�=��YW�	tӁ(l��]C�0�f:�R+62��	�y����u����j��{D�Jd���Q���5Jl�wTm���okc��5�jC�lV�r�{0y_��J�_�w\$�d�bhS`�	T�#^��1={�"=���"L���?�#CV]MY����a���Yl���$�u�Vb��XN��V��T)W�N����I̤7�3�Z=��}�p7�R��~��ʚ���=��~�4�c�EZ��0��:���]����Q;�[��z�j1�{���)U-�a�D�G�N�S����r���J0s�N<��K+�9)���"�˿�Q�j�z,Te��1��%>�;���&�)X%	w��:j�yh��勤v_C�$�Q����OJ��|5w�L>�_�C��� � %Y����V� ccv� ����(L;b����D9��<G�ƨ^���
m�Ŀ�V�~��`�1Ϛ���L p��W�+�^[��r�?(�N���dX��B.-V��?�Y���,[��%��h����bO�������ǟ��pA���oy��� BGu	�g�Sqns5_���q��U}�S<����G��
�M4�؊F �Z��o7�y�>!ާ���,�gy%��]%�ɷ�����nk��q���z�=���wex̲@X��{��HA��F�u��Խ�),�6�،�Ѯ��<�EG�tԂ.����2�x�"����^#�4�$�U��u!�_êA���$[��[�?�j������!_�ɾ3���v��Z �j=U	�e0ޟa��R+ێ�	�Ѣ��t@����n�?zn���:�z��y	�J'�+}��}#��'L� �r��c�$r�3׀������eG���?"�"zL_S��֡��P�|����b����ݿ�p?4vgq+/2�q�P{��� �B#�Nǣ�w�:=g��k�1H`gO26�����,0�5�>`�΃[cYˤ��tN�TY~h� �{n_D�M�F��쨿��>�$C*�ca=1�;� >t��܏ڧ3��l+��=�uR�z�笖�Gs��y�L�@�Ä/��>P:֫n����AE~پ�����N�����i1�����7�w�|:&�6��6'�1�gYt��W��Eՙ[as���v}YԬ���Z���[T!?u�'�؁~�Q
��e#��F�C�U.�w�Y���4$�A~���7�JR�w��6P݌f��ޚt0�Λ)��UԠK�ZF'F�+�/**����*��W=���*��F1�^��l�YC�+?S
 �N	(�J{iN�Zz��ߏL7#=e��(��Qn��޾�Aѣcm��'&$e�z�TI	�}P�dҬA:d��0?�݇<#�-��3u�F�b�~����y}�Ѣ�`���=�EU^Go����N3�c)�pdvQΘ��Q/K�$ETS�$i.9��3�fsB �n��팩}D�HA$��K:Z_�[P�p��>t�I���p���s�@Z�p`=@vah1<���Jہ�c ,qvZ�D�Z!�2������.�?d�{�趌i��\C���J�\�~�?��C�6#e��q�	w��y���1�C��k$�!<�r�>@&�	m���tfp���mܨ����b��>M��O��W��O�M�Z�>�Y�YK��l�(���qm�q�"RoTb�]i�`��W�4G�/����� &z�e�G�_'(20l9��#�����^L�`#�H���<� ,X�&�3��D���X0��- O;"�lB�5D��h;�fR��-��QN6�}2T?@	GP"�6��۰(^"�o��1�'G̫g�/���ѵW�Rg�=Ӣ���Җ�u�>ȼO��`K���Lj2+�q{�_?f�2�+��e%���a2�|���q�:Y�dc��}g(J6��Vչ>ɚÞ���lU:}��Y��V(}m�����A#lC�O�J��sc��d�������ǳIW�v�����j%b'~�}�S�P���[\�MF����OL;5��8��B-�{f�%̦T�����B���U�y6Hm�%#�°YP�V���yR�%�ʹ�k㢳��cЭs�� ��m4V���t=�� ����"��V�BGĚaA�)�ʟ��%���w�{�� �<��{2�˰ʳ���_E��DeC��<�1K:��wX`��tK���{�l���1]�4�K9�N��zij����ɡ
Vg��BB�H:���Ó;<.<4��d��!�]V��[jv>H�q���;}1.�pg�nφE��a�x�p_������v��/��d� X`��<T��*�RI������ʰ��t �f%�3���o=F"1-�ɋ��'Y+���a�J�&	H -���x%-Y����s�"�Pd��Rp��Y�W��/v��_2Y�Z�8�[$n+���˛���yA���L����le���4"n����?�z�@���+z�L��v���5��\��9��k�f�50N�r<�&Z=��dP{�6�ׁ7�����0�p���;�3�~	�P�aՏo#�>�b$�s�b��z�rzM�ky���N��X�Fo[ �(V8�ĒiI�Y��Ȕ�n�=j&3��O1��[
��X�`�ڍB���eX ����9�'��`�w< �����j�t�yy��4��-f#�x�L����1�t�f�|�6�P'���5��,����}~&I�h8��m��mc6?��U���a7䉀��8u[�$;K1v?a
����o6���-w�*�M��	��6��}���S�Q��j����<C����X���}O��N����m����L���F|�:�T�ߢ�=��<�7�
(I��W��+〒��I��r�����v��d7t�.$(����� ��Y�y�;k/q�?|����y=OM��El1Aq����5Ҩ�I����Y�j <�ϡg�Ǿ��N�Dw�ï``����i�S����2),�T� T����N;��q��|JA��ZY���lk*�DŢ�)/��)X�DFc%X|_ҕ���;��&���J9�	PLԲe�����!d(�\4[����~
O���$����h��* �^�p��},�7�ſ��#��</�N�t��愦ڂ�W� 4�e�!�4�R�CA��.��;���M�_X{�=w�*��#�3@���k��7X�#�gfn�Ų��
�9��QT�LEP�����R�@$���qr	
�BJȰ!�w��#�mx����s��R�:26�JТ�o�]���b��:�%�`b���z�Q{�R�0QB�J�l{�ɐ��S$Qy�>%nYkR��8xc��7=d����TbٵQ0ޙ��}��r2�:`�!�B��z�>�6h`��փx�,<4 �O{BVA@Q�Q���Et���XtмF���iOQ�?��U�n�`��q��Y��L!�0�]���� �p��ZFX�zr��7���,'����U�(�~56<Z��HL�3@�����D�eZ�7��!��4:�(K ]��MF~��סr�gxߗ[e�M*@�W�
I��*�`�����.0za]���6>������/`�z�kQ۳�lSu�s4>U������٢.NbV�$r�e�X\w�� �M\�>�� xP��À�/��V�/�c���31@��%1L��D6�1�C��W�`7���].��i$N:���C�׬ψ=��L�E�M�*��[�����܎�K*`�<֘�$���n���[�)���K��h�F/�	U<!q�Oy�\9��	L�I�{���6j�� v�gVA�����;TS㸪��V?d�������T4*�0wt�$��ۣԖ��u�+��L4DBе?�p��0���'�~��%��l|x�ڒ@�P��&����s�����ا����ߊ��C��)D`\	աVd�����}<
|�]xC�NuI[����2������<F��P�7�$rl��A���*��A��W��θ���݋��`����E<�rP���(�d0�'���O�p�~��M�M�������~C�'�f�]� :<o�t�P�gO���6v�)�/���Қ�e�\I���t�$9L������w�e3���n+�$�U�*��1�r�/ڕ���������Pj�"��/b:`OC4�Z�����${�~��Ź�?�S+��h�-�tF8J %�Ny%w����˯�+�F"4��]��>X�c�A_Sp��o�E��!���u�M��t���߲�T^ڣؽ�G4,��al\[��z6H��6���ʆ�X�}����p��P��\���{�]��ؘ���[m�C?�	@��`-Q�V��+!����4Q����T��V��f5BFc&e��;y
?+�������~��	)�����u��C9���F9�F�7q&r�Y)�����}���N�'כ�R~�uI�Q���Nd��Ք[������i?�� 02�l&�F�TK3&
���i(w[�6)P�meQ[�/='v�B� ���Ξ���fk�{�&L�l"��撿0A�W[({����������^b!M��p7|tm���̺�܊��:\��b�&=
����Uxk�)��Ńг�4�Q�.	�\��K$k��n���.���K�3�,��r�(�/����1��Az]Q"�� ����ͯ�S03|�cX��6
Ć>G�+����3�� 5��
�I������bp��|ʓkF�J��*�&�����e/��I��ݻ��V�g���ĥL1V�W��
c�������5/�CuΛ|�]?��8@4���o�[\�2lPA�<d&�<{�i�Vo��+����%9�4�iO�=9��kS44���&���W��}5�_��FM�-{ǒ�d�b;�_�B{��!�fT�|��n�p���d�vG���oǇ�'{5t����D��bw��m�����A�7iγѝ�Z�6nf]&�=����@��p�sߩ��4��^!J*�֐To5�c�r$#o$�ɧ��F��E��jwu��F�S�?���b�v�N�y��{����q�L������`��X� j˹����6*s�����9�!��nNɌw�o=Al�� ��S�b&�̐�~�r6��t�{F��&֍qc�T1Z ]*C�Zi�fkn�a�T �M��H)`�vn�>P"rs������&������6?�����T�ҍ�$��VTP�{�T��1�L�����#yl챕��	�� �n�R϶�l=�
'��M���p<Ԭ���}cw^�^@aOc�af�����4�|��iv#�_2����3�2�K��od���3��]�����z	\Qp" ���#�!�F����F���1�qzWf��Tx�z�)���6���&�j@&�HK��Ϻ��.'^�T^۵������0�m5<��a�߀�W�O��zN�0Y��D ���ę˿��N!ÁL�����F(�������k�0H��Yb�JӠCfj�S
WX��-���m�o�=O�KwҔ|Q"F�@l;hʶ�XF@n0�=��XH�h@�K�Pš`�σ� ����Rsr��Pq���8$$c�Z�Es�fl�����mD+���6QN��D�F�o�m�;��{A �nM��8� %����9�5�Y^|�X}6�Q������(;��E�y���CIR�?�U_�U)�Hr�S�o�^]��U��}�{l���`/����e+O+߯�_�΍��1h�d�&�KϣK=)����1�ϖɜ�r8�����͘�v9�7{c�5�s�>l?!V����Zx��R[���Vn���MO#�t�t� �#��f��m#MY~c�H8����п�=�N��š��}��}*B�t@���X��Je��<:�sЂ��V�u>fP3֟e���#�zdu]*c���y%�<š��7�V�w�� ��a��v�hX��+cc
�:SX���O�9x8u-l��������j��s���ׅ?��v7;rU����-�_�4��Z��|�z�~`'��X	����+%�����Sl�5v76#W�<����{=�6��cfK��/�Z2b�WK)*=��.|�*� Jp�)������\8��A�m���N�/�*�5� 8��e.+�������y��c�2	�t��'T���L�n_h ���q�րn+�]�(f<�P%�&�h�3 �̬���h���閻�P��q,�}�_]�.(��~�V|��L��9/��B[��	Zo�Z�'%�z rb�뜍��'uQ������U��X��u&"#�D[�e����x��\Si׬[�y��L�/�M����+�T1-�m#�2gy�ry�7C�~1C(K2��&��Avė����~\4I�J ��ן^�:/#=@)_I�6���ɒ���UUfY�!�^}y|�i��a71ʾ�I,@^��-�k���qӤ4��:�dbu�9�` m`�!�e�W�'�N���碉V����'���`��Y�{
k�vT�x'JzH��I���?ow6�P�ƜYK5�^�q2����z~<z=(�de"Q��B����XHM�i6`��(~9x,S<2 ����>���B�ڬ,K�c����zwGW���EĊ}%�a��0�
�]�������v^��dl�[����+�Z:^&�[!C2�?Ui�\ᦍ�oi�#x���Bho_��Hð�\�}�����@�K���N˅���i=�{�"{���:�Y~-��fe����@Zb�`��.�4r�`����Vu�D��Ջ
Iߒ+ø[�������*�rg����A� �⡓��v�<`�{	|��V7ށ�k��	ƳX�-s�>��y4�a�<�K!�+c[}�U/0_�p����
�*�I��_�T�Y�W�
̴���%$�`w��sS��
�ֳ�#�
Y��=g��?\��6y�*Nϒ�%E�_�l�Y J���(�|��k���/�?e�&����T�mk��脽e�d��{#
�����w�=�Q�'�a�j	��f��Z����462{�*i����tm����Pi�[pBW�u'V���Ln�V�Oo�Qt��eX����l~��}@��iۂ(Xd��VW_�r�ce��3����{����]&2�T2�o���'��5�F�Ii����5y�F�ƣ(U�������!�q�� ���E�SX�ԓ�AzmZ��K����[���9�+d/NJ#���J�b����بɩw[�#��$���:뚿 ?��q�^�X�$����N�2��/�*ɴ�<"N�9uֺt�d3ܺ�b\�Y_$���u�\JtP;ZBn�t�K4�l��-NڵGil��D���P��&��sp�"����B�T���i�v5��	�w�K���᭖�4/j�,�?}/O����ש�M3�K�M�`�|թer�A�3��62���n�kI�%Z?�f��4�	jR�
������t.I!j[9z�G�>ՑwS�M����}h�/����u
�9�#H�E�ha	������zO���1���ί0�!�"��ڳ���A<F�*E��[��Iu r`΅;�]k���@�(�i�R�T4� ���i�C�S�M�Sc���jL����Y �ó��\ڏ�FT ӡ��	W��\`��냞��a�f� 7M�������H YR�I��8/^=����bܒI������H�5�0�Y������r�F�ٜ"��Rq�_����[�+Υ��x�Vx{���B�Wb�/=�3$DY�ɫ�Db����d��b�\e���G�$���s�<�9�|P�GH�H~2���]d�k�c�Ø�*�i�х4MPxE�0C�j��dr%�<X����g�D�n�F�Z�
�؍n��,2��6u�0�Y�='�ۂE.��_);�U�D���Q�aa���zG���|�#�;����Ę��`����E���W�D�p�r��� ���Т���EC,��&�\��꭭S�B�������4[d��|đ�Z[�2�u�x,�/^��x֢I��:WD�f�74�b���Ǐ_����5��ay���d�%�X�7�쌠X���&�!.�XCn0�����ם����e?ڙ��=�u7'�5F[���z3J�'��9�$�/c�}�rEE������&�fŐ�)L��P�;y(&�c��l4.Iy��`�G%By)�i��L�Wk�lu�f��Ŏ[�殟/Քܔ�O��a����m�!X��|,�=�=p�S^��0m�߹�-�sj3b~JF�/�nw`�o�w�\DkR1��2�ǳ&���V�j��:|�P�o�����(\��:\��?3,%p�ߎ9�����VY��³�m��[�J�K���m�:�)�W�-�
Z�frN�Ś�SI�N[�:��4�ȅ��b����.�a�"������t<G�{G��E��a ~[�/8�'��<S�j�`
	���+�Ä/�����X����)f�R,�ix���֐]�7�*ט�$�.g�~
��Cy�s�>-�3���B������A�!2 �=��́~`������
N��P��&h:�v��� Ϊ󏇢䌥"�Ͻ�_ɸ"��j6 U���̌W�Z�;F�$�DEa�aD�{�����WnIGI�Ŀ�Q
�<P<�\�,5_�]KG�9�F�"T�������5�2��cN��吃��a���~�ؓ�� .��kM<Z�vC����@��2\aYLI|(��o�Q�C_UʯT��ǬE��;ê�?��оZ�89��@� �E��e1�a3�q^]�H�5��S���I�H�jgh�
���ؤ�'aDr��1夬>�TN跢P4&B��P���.�������ԗ���<��Jbذ@蕱����>A���X�7���M�X��Go��� <HP��e]����"�l�cׅ��4�H�Z-����"Z(����7��q�B��9u�TDeѺ� mΨ33�,�h��*�O�1��#v_Ϻ�����WZ2��&yPyI���������a��l���n��\;3>¡=�qgܵ�� ^����qe�,I+�U��2���1}k����_'�N��M�OI?�~��W@`,���亶?�L_?�*9$�W7e���� �v�`�FRL_*�����Q����d}�����{ 9��w��2��I)�������˃���5�y�j��pP��8�<��h�q	8��D��݇D4�L�Z���򫎖�|h+�H}s��{A>�
�@?��"��UZ��orq���ִAr%��f��Y�2,��X����^q'�گ>��}s�� #��?͗7�;�˝�@�i�]��V�gn���EӜbj���ž�Og'� ������ܘ��׎u!�9H���)�yB��D���Q��{�`L<����͋����N�T�:/~=i��a�������mdҗ��.F�&k��F`�jhF�o��A��|Z����A�0��V��仗Z�Q��ݿZ��9x�&�r����W��V^
�mW��p�4C�iM���|�Ŋ��(�h]�4�ɥ�Um)�N *��]g��ζ���Ѹ����9��50)0�st �4��8�]��K����+D̿Tw�`'�I*�ͭ�El��FlA�F7�� 1n*@,a�ox�g�!��	��q����B�h^Z~?t�"�$����r���A=�ȍo��L��|Ѝ���vuJ�N��(��.j���~ǜh����M����X�느��|�+���P0Q]���"�|6�_KO�)�����l���e�7�p��<�{�	e�/IFݰ�Gʁ���]sr�tZ����	9��Ta����@����R0�"�Ku��$T��ҳ��`z]}L@l,�+h�C���5"	�mx$@�\�Ms`�q� ����Gl�;��CKO���F���Y�!�y�jr�D���⭓_<۸�OEd��r�����B�=)��q{9���V�Q�3�K�������i5%��1���~@�ئ�s]�p��p.���t�RGUW�Q��'}0�ӛA�-���]��cN�Z��&Hb#䇋��Ge�(���|!<�9�c��3��{i���*���R�jK�� b��0�(�;_�I���^m�;>r�S�usM!�6E����f������f�S]��҃Ǩ|��*�~<%f_�Ȼ���&b -C�Ɂƭ![;o>���m{��I2��T-�2�~��P�-y0�iH*Ƈy��e.F��Hk3Gu�����#��XK�Oz��w܈�\���і��%�ie�����s�̓��q7g�C4ؠ��c��ЎL-�F��F/θ神XW&՟�MJ��_rR�6 ex��^�����b�%���ѽ�Jȵx��0LPV�%Y��m){W�п
���@"{6H�K�&.t�z6�8<~����Bi�l�����z��M�X��K��Ug�_Kn^��8
i�żtf���єf��
�>��}䁯#�عN�'帊�� pH/��0�em��n�"3k�6�$j��\@W�>k�]�^�8�ȻY"fX�G��$'=<:`#��e	
�NJ*ME0�֋��t��1�4�b��>�>L�H���<O��Ϡ�������W�Zly�dlrow�ᦛ���Z1�Ra����4)��l!�3����AX��~��g�W�o<|���K�a�4��A.���}؏�
�,	&^A�pŞ�0l2*�_��
�B��_�����jO��5f��<��Kʋ�J�X�M�C�y��4��"ģ�iK�2�o�o����X:H���v9ۥi١��p27��zS<T���f�˦q��������M蔶��Y��[1�3>��KD��aD����W2 �Ӱ�s9�K�DV�|�w[��*~��tN	��D8��k��nh֋З���N3��!���-r��_Bz�5{4�fw,�w�[��Q�ME�lka�E�6���zC ʶiq�x����%ˉ$~�L�8N�Vݷ)s*ee�7^n���S�abs�T�v������P�q׉����F��`	�\�\}���b��c?��h~$5��9�P�7��m��-T���k��殂u�Ϧv�t�%�X��Ȥ�5щ��BƓ̨��9�B�Xꈊ�$,%�*�ire�~iy��R�i&��Rt^5Ù*�!�5���1#e�f-���B�c���ҷ�u�9�����dHs�F�[�|�΋#<U;��V�fb����y�˰0�T7u��1�}B9G�tٺ�p��!,�m�=�#�	�/숷gv�d�H��.EP�h=iA2�'�c#u�b�	1�.�I�ZA���.�kʃ;8���z��l��]Gl>Y2sxV���b�oa� B=�?4��Ҍ����#u^�����y�a��fN3��𨯆���x+��g�*el,��V�v)�v;i_"eb�d#�\,'S0�bf��#h�K�甧G��. g"�Dg�v���b{�L�&l�
�u��g���)3��jM>���駒d؊�p�MO)�d�y��F��%�[�����Hx��ftR]��Mْ�n����qZ�����[Qng(�@�{�����a�[.��ؑ@w.�$��J��ʑ�n.���R���
�ϩ�s�Vi���c�9�U4Ч0b;%5f�)���t>��B��@��Xp.���,G�����H������_<e9��oW�c1N���D"޸s����-�H�(0B�%ç�R"�<�V�MaF�H�9��Cd��3��T'�<[i�[�z.��=�'��*ᖊ�)�u�Hz�n�ڗ���msh'Ľۭ�^p��ƤOp^\"3fC�d3EH#���Aw�_�.{�ӳ3�V�r���􊹓>f��[�Ƙ���f����*	`��^��r���y
�|(Q�С��.����`?K#�P�"�.���7��"%����x���3<!��]�!ws��wwN��5xU������R�p��L.'�0X�;��׽�p����������=Zm=C�Wݭ�%��jB�	�>�f�1�W�4h��cQ�Sd?٨A���K�މ����ZaÞ�Q]) �2�xN�����] >S����'	�uMZk�#5$ =�Vcq9��\NŧRB���k�D��PBz��$ce��4�.����
`�pEJI�YQ���E��{���h��u5?��G"n�*k�J6���'�ü���na��ȫ��3���Ju�{+d��"̑���]l���NP/���.������m�D"�P7���$�r�C�7�����vP�D�٫�8���m�J�H�3���1Y0�odz��&��x۵�7;�lɁKV�uhf"j(i@
��n���*�K)��@�\w�pG-mD�<�Vf�j�x��)Y9c6��``�oW;������3�����T5 ��h���M8�� $q<u!�OP���0������K�;T;5ұ���-���3h⪘��ގV%�w;��r��RɅ6V�D��y��o�n����`<�Ns~�:v�[q��Ѝ��2n5���R�R�wk�YЦ��	'w��b��2�5-�P�'�l@�8i��T����v��YA����C8��ǿ�&�u�Zu
Յ�j�ɸ��W~?�{&6�S���4<�s(��,�t�F؋~��r�9��7u�-)�E�h�K���Oi��1�켕!�M����Sz�)g,QFC-�QDI��+���%|)�_�4�|��EY��Յl��O�`,���Mq��s�u�"
|ǣX�͚��B�t����rmt�,��7a'ȕ��N�'��9'�_��z��-�6��4��:�eo�����օ�o�r�oޚ��Q)�A�$��qG�)1��t{��}c�rW �$�g�ȞZ��E���Ҡ� %<^���[R�R�F��g�j��y���&uZ��!.��>��'V@���kʱȠ˲��*�1�S���NZ�$�I�mJ��u���+�����sW@��{	rŖ��N@���TY9��k���+�D%`�;�
ʠ�[�^Uy���:e�p�<Cz�yQ��ȳT �>�g1�{�s([R���y����mT/�:F��8eI�|�3X~w����8�iz�y9)���X����å^\�`���7������'�͓�+f4twٟΘ������E��0���s�$t�?t�3�I�f��S���2či����d5��o�eGV>����O2��mh������qԍ�9�4,Ԝ��7����}����+��F��^��ޡ
|��F��fSZ�,��>��.
�K�ࡆwC|�!Vw-!�$��eV�ݾsY�5��s�_�x��S���\�
,�؄'Eox-DM!V��?���|��4XV���-k�lp^�_�����E�������3q�?�TK���%\�ݒ�R��������K��[��5 C9n�����W���ˌ�B�ܯ�$����J�V�@�)� %s%�MG���ghO�~���J6;z�:1�bŕ.��;YxŪJ� '�B�F����zl.�S7��$P�/=ɲ�3%�]���I��y�#��	�^�'	]���<�p�O�3.�1�y$��٨�7������{_�5�Q;�7����Eꟻ��uw~I PL?q��řY��F�����Q��eu�y�,����0�����u����E����?\\��`��Fh'迻��"ᱳ�!&�
S�=��3�X԰��L�{�5l2N]�$%@E�z�J�WN����4��@U��D�(d�{�A??�t�I���蘋~�����1�SC�	r�>�U��i �5O0F��X�[��{���N�"�^J/���lہ�H5��z����?�6J&x�f�Ǝ`�5��7?�T3m��@��+t_�|�-\y��o,����H���#�$U?�I�)�%bn�k�5���o��N$#I��/�����(��V�?��
;,�AH|����oP',W�� �&���aM�q�e.=8���G-����ӆ��D���7�#�#4��ˤ��-*��/6�r�&.�0���_��j_dѱD��ӳ�Aj�?2��Lb�P���^h�2e�t�@�L��<}Z��`&&�~!Ĥ���s`q
&A�5Ae�J��Ձ���I�� �۳;u���D��\M_1|ה��i\9�bT����.@�Qe��-Z;vr풿� �����Χ�:��a��l
N���Z':���/hOj>��k٬�Q���54euɁ����sr��F��5P1EMuDtoR��	���Ik4���%$��(��U��٥w��e���>_v��]q�g䌊�4���Ўx�C��Z��O�}�E�~Pf�;����yK�/,�[���I^����M{���~%�˴\��S��G͢��/)}\�m2"�=���Ԑ9W-[��f���ҹk����̖3ԯ=p���Gwq;��[�+���k?h˕��9xv	�Q�������͙G3���1��jv��Y(��)�\����*�n�w��&�f���[�(��e{q���]��uwsU*GpO�S02hrmj�G�5	6*T��҆�Ȝ�d�?#/�4H�r�����Z�������?^1�18S`M��l���S�q&�0~�. *�X��<�z��:J�'ƪ����
�P�[��j�
����G�#�q_���J��ˑ�~q+ �N1��?�(kN�Qt��gw�_���1���ϧq`3u���q��_�I�i/ۍ'�C���8n>,��ر}>()�K�<�_�����������p9R�
ItBK@f��|�V e{߿�&3����4�i1rZ4:�� ��N�~2~��U��EZ��C��N�~�̦s�j��(������x��0�=���.�I�͚���R�k=e�/]Rr6#�W�����s��yQa�h�)ۮ֧c)��D!}K���KN>��8��id�n�:*E&&'zrv&���E6d�eCu�!��)���tMV(٣ͽ��*�V8Cj�+5R��(y����y�cѹ+�!�T�O�
i��3D�D�Pќqa�p5{���v��|���0f�B��{t�|W Rt���� >��:��n��]�c�'�T|EKE9<e�ɑ:���j��wu��C�VH�|�2�U�y*���� -�&����i���O��i?���j������4D�����u�u`t��NF�[���&U�o|x8���}W�v�]D�0��� �̪?ր[�TnX3��$��$��i����3��<�x݆*G*z=]��'-�c!C����'FX3�D�Fۭ�F�Jb��g��� �
^���KL�λ��gn�f��?G�H���໧��V�(�lG�_G�|)��zAN�O���WoM���'��t��͠�4��W�AA��h�|�t�RA}�cNr�g�c��� C�N�F$[�v�<9l�d��5�g�B ��W���Y�ġ�(R�ռ��q ���9�H͞���Vv^#G�y<�2��)�l�H�;F��}'S3�
��� �X����JJI�ߧg�,�
'i>dU�v�-�j���j���y*! ���m�0dU_�j����d�G��Y�3�ypg�D�)�����c����C|��*�}�����XZ�aq����N+����/���IbL�C-%\q#�9��Ⅾ�����g��A��᫠4��K��bNm!���sN^�Z��1=�:��P	J���x��b����w"vPH�)o�L����ɘ�n$k�e�ͭ���y�`	�"��#$��h�5�3�3��d��V�(R��G/���?�}{�"�O��*tª[�o�$�ڕ�$vy\\���]�t��;pxh:���E�8KnxZ�,�YX���a���8vŨ&"�S����wɺB�q�q��:��&'�O ;�4�Ƿ�'��Y���"�`l#_EȦ$�j��AR�V, KD������rnj���_��d�ց��
���X1���PN�J�c9f�ȧ�#�]�VZ��PJ���Rx��Iz�hXs����gG��3J��?���`�(���B�#����q�<G�$��W.|����+&��7�:)ǟz�Dc[����ٺ�9��*�~�(�įQ�**P����־n�'1A��6�#��2JX��S�Ɣ���g��ot̹8���
�jy��Ʃ�|;��w�Q��]��C*v�P�,�@�v�<�����|v�mc�d���������k�\+[���]�xd�u��M+���S|+f���^\�����5�G��W����L���jE�N��b
&�=R�h�gq�@^���]������Nb���ʙ�8�1@��� CcL���nEk�Cq�1����~,�4�
���;�jW6&�]$	��q�Q����K7*W��G��y�
��;*cN�]���B�N+�^��wK�$������Sc1�6Q.6}^�H�Ѫ(�1�ի*.�+�Y��׀Q1X0���o���})�Z9�{�e���� ;��JggR��.�*f6,f=Q��l�r�;�$�އ����ɾ�!�����9\�ZR'�)�Noӡ�v_�0?����7����BG�/O�4F�fpx,�E����v��P��j
¸���2���pa�%���B_?P�y�����u��?��i8��F��AR���B��0v�jQ��t����O?G��0O����MLw2�j��qwR�FB��T7�5גeܯA�`����έg��՘/M6��!�f�Q,��ϲTo͑��1�y��-A�̂ ���ݽ�s� ��N�Y�T�`��XF��(V���D�<�vf>����8;sjm�c�~Аj��/�z��g�K'��BA�q�t���3�^��	Jn�4y�bj~�A	��9��u{w�\̅F$��wvs!�ViT��ˀ���i�!�E⼺ �T��I�viģg�Rek|�p'=Bp0B=�Q���p��4Bj[�3�^���r���>	i��|܇E�Qg<nZU�K�����zȦm�ZI��8��ơc` ǰǮ��U+����c����Ôd�p� �Zv��*m*-�n�E�A>"8*�V��:�O�tJ�H��r�b�V�����k�LY~�hr%��H�b����5��*EE�1��3�!S��#c���- +5�5�7���edYXJ�Ta��c�6?�|m�F�9�����a��Q2�������1���'��쎙�JLZ!K�V�{��M=�?��K��`��q$rF���Z�w$�Uث3w�u�~j��q�������5_q�H�KLʔ���z��9�*HCW��)������ύ�M	@��\A�2}2MS|�[T�qR+<��2�&'�՝�C���kk���^�c
*�{�������=�(<��(+���a4�8���CԤ��5����ܩ!��D5ʏ�6��G��HW�o�S��3
;�)�T��h'S	�':�XN�&B�B]���gy�'��I1e;�U�fhg}��%�@���9<��&bsz�ϫ�/�sE�; ��iNH�;{�N=9(��z"��1���V�C}�,K�c�r�\�'�#��§�`u�K���մc���]Ilu����tW2�h�+L�^��p�a伜r7c�bD��w�˩j�Zvf��EW/#.�)Geg�5-�y
�k1d-�^
�k�`�z�
Y����z'4w�S��25pg~k�Fol<��}�e�, "؎���f��e<̏'�Ae�Ќ��r���P�ǉX��9��S$M��;L����Ϭ|�ϫ�g�����ŋ�
�Pw�=�o��;<ёf~�j��
��O�y����14�hO�ʔ��-�w8���^�ʹo��_`V�*�5ڜ[#1���EC���φ'�"��#�Q-�W�PD�F��7�Z����蒞���	����G�L���Q�iULF�-[���[{�f���ތ,��)��I(�_�&�"ws�|ZN�A�AX��
�G��Y��*��tp��R����T�>�؁�!ࡦ=}��VQ��[m@�,�!YΦ�����Ѐ���%��u�^ �y��� �Ax�]��Qs,�f��T^1�$�5I��,
%U��#�%e��NU�O�Fu��uvI}
�����{;��k��Ds�`����|)G{�:P���?��q+^م�]�XǬƧ�y��1r��=y�4�%��K��
|�n�pF[?ި���1K}�ؿi�2$�7#�VҞ�,��n�|�H���>�bV���l^�C^����5��j��
�-� IP��9���dJ���i!ʏ�N�1m��{y���PCH��H$lV4�k��5@8��{`��d�rYQ�kܠ:��:�@e\�� 3`g#���<��*ӡ�gg%a��ں$,	��&�N����N���i�
�GR{�I�{�Q�*���aϹ|�&_2w+Q�g��05w^C��͙���5�sl�퍧�'vhj��
0�9ѹ�	�m���_H���Y���U3XQ��+�c 1��\�ڄ �0!��9� ��*�y�H�kR7������nE��n����܍+@�9~�}��t�՝�8w��J���I��&5IY���
l�?=+T��k�����V�hH�կ4|���^�	�V���f-�Y}�i�4ɐ�����]~����)8���_Qi'>1s �S�IBj�}Ѧ��5/|�s�o�@�ֻ����-����/^�~UG��_��G�\I�ci��(���6��TxV�y�3���e~+�F�V���d�P��)l�Q0V�)9�`\��Lɱb1T��i�������<ѧ`�O�/��o����4G]\kmR߭��~����Kn��[�ϱ?koE�����7,���$�'O�(��u�/��x���8��6��pX�W���<�hw���G�~�>��c_��m:�)~���v.b�5\�,H�1'��\Q�om���]��
4T��Y@�W��l��Sp*39��V�`3�	�n�swf��;C���o����hJ������ʋ�pM�)��-a�E����VMɦ?rƁ�h�V~���(0y��$-;�nh+2�`<ْ��"u�CH �����ȝ�v5iE�����h���Z�k	�4-�[�'�t3��t-m��Vu���f��qmT�O�4��I�T�w*�c*Ŝ@���P1�(��]H�I��#Dz���JN��]~��*�EE_8���]�����,��^<BlC�a&��M̯f�8|CnzE�h�p��y�C������w�.Dy#�5o��p�*)�/�PS߄6G´J���E����$K��Gh*�r��we5F
whs=�+;�g\p�����#�!"+'���[Ŀ�|�)AʾҒ��Tv��C��;߇j�W;T��4��]�Y1��;	�UN>Nľ��"��g���[[���4�q�D�J� E���7Q��g�b�c]�͝~B��-u���P_�\�U���E�%^���j
�tO��)"��k���R����0Wf�J�AA	��>S�8�\���%!��{�҅���\�ae֩��ܟv+�`�:p/99Tڢ�h��R��7 ��qe�E�?�E��rrr�oL�n:�L	�G_jD�>���N��E���׻،�D�8�g�	���vH컼)H�pΙy�̀�	�䚮z�e����`X9�<������{'��� ���'k�)���ʷ����b�_�G������cNm��Z� ��J�!qiK��Q �����s,��c�3ojz����O�?�1=`��:~�k�ja�; �5c{�z��f��� �s�Me]�ta*#)R�]�[=�F�<;�0H@ў�(si�}�����bFA�W�̀�y���@�z�(�����F�fvz��i��?o�B2��7h+џ/��F)��|�ي�m����q-[h��/>�Nh����2v�E-�q�ɬ����kcZ�ގ>���ԃ���9G��.ET��O1Z�hf�z?�/��W�'�$����e(噔��cs������@_��ʜH@u��K6c7_��VW��?*{ku@.�p-�{���"���(���K*���	t>��<? �N�&�<�ɇ�m�g��������_�<Wź<Udf^<�$�4U�0�~���]�~Q%�>
�e�t��3�ı��$��tgG�1��P�R�Do%�2g8�~�m���V�P�����ѤH n����5Ť~�^8[`�_!-n�V� ���w�Ӻ��"��{|�ı;�V��1r�O����gD�3�J��
�ne�:3��I���!�2���h��6��dnLGW:�\C�<O@�k{���rg!�ܶ�(=�42�̀y��X������5Y�����!:e �|f�u�z~YaG��l�����%z���}������I�ґ�&e��P�J��O�|��K��*��'^%�2�';�^>�n�I#�RF��~k�xd�O�ܨ�M����z�d�ӝ�f:�=��`U���@���YvG���/f�ll$����^��E�fOF�h�����QP0�;f����@�`��bb<�\���V���*���&��-v4�Cg�T�:ZE�e0�h����<f����u�������5�� Ly�~���� �C�d����z������چ�w�Z㰍�v����חf��89�"
@���v�i��گ'��/;�fv��󯫦��hոy���{Y��ߏ�x����p��I��/��W}��m3��O�.&�x �\�����V�`NR�4�&�]/�Zw�4�Ú��~<�t���Q���i�Z0�4o�w"J��+N��E('b6W�2H��������ayY���Ҕ(u��tZJ�yb�_� ��EW}󾱭Pf�Ʃ/^\ʮ=�]ՍlD�����,We@���O�G�[`�	x��П-#J&=D�}N'bR�y�v�E)Ó � wT?�i��z��d�B'9�T�d[rlٮ)ֵPg��1Wp�z�榟 ��
�$��8t�ΐ�"BeYV��׽���7�C|	�ܐ�]���x���BV5��6�T�
�-�N��/i@D�?���b�/k2�'��h,�B{2�D�n7��Mڋ�:��y<@N�R��J�*L��0�-�jJ�ͭbv��-��<qe+R��r�]�Я��J�e����ך��g�� Y�ddו��A�e,�G?��}f�,Ũ���;1��lz��G��s�������,1r�`�Q����
͙��6��"R@�} ܲ�i1�}��q]o����De2]�ܩ�j��u�3��v�bL�8b�)��ȕ�N�'���{E��i%������F��Y,�a
���@���5���s'p��le�({M����K~|�mvLu��0h�tv������睡�b!�w�D�!�ΣNz.{*�H�3f�ɬ],��_l�s�E��ߔY2�N㻟�KO ��`l.U�Zt�DGY�m�c���0�lw�(��ɜ?�N����-�]��_�;��S#l��9�b ���
��ɀi���=�Ë��>Qz�H�^4P_wL��"%'i��yg�'.)azn�6{?k�x�񠺽B��*Ĺ:ȇ�\g�񲬶\U�EJ��&��Į0a9Ȏ�Ʈ��ޡ!�%���}��������`œ�/�jG+�j�!�k�����Ӏ�0dQUP�98������U�H",���%��1Q�k�d��%�����43�>Ÿ-���R斾j��t�����f�6�pm�XI�Ae�t!�M��UtM�U�;j�PY2�"�v҉*��#���>jy1K#�\�'�dky�
2�)Dah3���,��/��V��؞KQM��$N�VL>�T`TU'�]��z9�K�$��N=B�N��\�Yq��.6
�]��a���f�|�~Ac��Ϝ|�׸�4U�H��z��m��)�eKՂ��dn�����E�<�$��.MҊk�yZj�N"C"�kO��&d�A7���e#��.�x�l�i��ΩY?4Z~H�E���W���1��T�/1���0�0�ڥ �j�K �&s�ۢLy�Hw��Z\��I~km��̿�hq,rϡ��Q?	����/]��l6�����׉�HYTh|���Z'  �z���T/f�s� ���jh\�%!�_|�Nʦɸ^(bJNm��+_�T&��,Pve��p�|{Gh���2�� Am��>�8㍢f����g'��$p�y�s�B�c��>'.J"*A�rɥ?�`��M]�&�
,�.V',�E�m�VI ��v�W�߭d��j]�|Ev�:�3zz?s@�uv[�d/rs;ŨK��w��MQ���G���7A�֕d�R4����Rfa����cwy�d�s�qo����q&{� ���ՎPd�Z<�
�n�YT(���gN�:��hAյ�3t�y�u~�A�-�7�2�^��9�=�Ie�&�4Sef2&$��.�:�N�I�R��K~�(%d7`Ʀ���rd������� �ZC�.z*��#�u
�XQ�f��ƜT�&������Y0��e0*@aw�r	cx����)�X=�>ś0��׫e�3���Z��^�Ҟ���2F���=2'y�SI7�����~�����L:'QAm�8�35��r���-����K;�$l��>�r��1�-ʂ���lg�MjL�߉2�b���@���@��E޸br�A�zu۶�/�8Ԓ�:���g�N�p,�R����&�2�aDք��oѰ�����V��U�W1�֜�3�a�=fq�?��XM�K��+�P��յ�f�
���v^(�n�w`C���gjjV���p�]i	�5KQ�LfVx��G.��,�Q5hȷ����IE�*S�(���v�d�t��kaP}8�Q��X������1%n�a��n,�oUN`AC�B�?���_`���*Ί
���;ƨ�qD�vCZ3
����xA�N��L!��u�)��#$=���/�B���Ze�n��z_�`��Vv򟏓P��UH���ץұɆ�z&��͇̖���D�3J>���I=p�*Na��
إ�C�b��w~���4�s �.)�|Pg0���
��n�ڟ����bZ�Pe�X� ���\~Z�|���c����T��8�>Å?f�zԏg\ZQ��o\�j~�^jS3IlN�Iz�h�@��~.&>n{�MBV>>!D�ܖE�z�{y�G�1��=��:a�ڻ���Q���d��i��]��D'�Ŕ�ZƋէE���s�k���F5��I&���TL�]��q�Fn���������}"�*"��Rnָ����E�~���&���?�ea<9N9���Ǿ!�Jz�gd�j�^%��4m���te�e�Ef?!&k�Q��r��e���m��.��7������E��Ք�a�r���k+�s|�QG!�;?l!(a�o��>G�Q����}�vI�7*o��B�$���h8�+�GF`FL����3�E'~v8Ns�c9a���6�V�[{y��]h�E|'���l
��J^��~�A�ˍi�p��1 Y��o����*�=�����|�32&-�]U�^+*.w%�a��z�]e���o��C��(�q2����ԅ��̈��2����d�K7�iMZ�a�v9��~ ��8<[0y͛�ڹ����:Vm���0�l0��c�,��Dw;�T�p�X%oz!��Q�I'F)m"�%j�N��=i����H�v�"Պ)� r&��[
E�Թ���](���U/]��9��̱g���mH�+��L�M�ᒉ���\8�ϡ�<oK>��z3�׫T���r}&��5�x&��N{d^��O&�9����^㛉 �v����j�v��"��x�'�Q5դ����u��r��^x!���:���qy��9�"w�\�{��H��	 n �+��moR�����ֲ94G1y�w�-�Z���]@!A��Г$��u���<,�ycۀ�ɋ2�	�vSt?�iYKZEB�/h�uV:���cE\�&�VY�\�z�Bvu��vx���A�&���Ԝ�8 E�\w�G���`k
#cu����4O��>��wE�-���2Ķ!���h��E��8���%j�F��N-��`z�+��zR)�Ƕ�r�q�ϯ��R�8Ѫi��<m,Y/�FVt�;w�*:������%����/�xꀞ>X���ˤ�U��}hY��ɩ�ڮ�L� ]��4�E+W��y�{���2���g�5�VP��v ��8YD��2���u^z,ΡjU���c�|�~]'�U��p�أs��$^Rw6Q\���A�1�z �E��|���^($׽�dv�0ec4 ��3��K.`�Wodn�{��+?��0��{2bھW�����#�fǇ
�k���NJ��GΏ��?�ا5��dIf��x��`B8�{�^���Ti�
��Ξ�sx����*���H1�߂8�@PN�� L�~�����eAG�H��I R�M� �p�ub^<�gǾ=�#\N��w[��f澋����Ms���4B�~�{b�q2p���s�Y�Y�����:&B��:�^�φ �����$���=��, ��m,h7$7��Ɏ5�hOu��{@��>��_\U�4A"~zn萼��j3�i-_?��ߛ�u�Q	�HC?���O�6R���+��5���^|�O�Nf��7�,�������2۸�]m��	�*@�^����P1���B����t�0JN��u$i�GKL����1���Ug}*�<]����rG�H�F΀�����M�%��vt�;�� �q���EN���/����]e�_�<܀���FդMz;#� �����_�9D�9��5�naG��sP�+���K��܈:kd����#R��y�������BDS�`�]�-؎��<�I~�\�<��x@Nd��?��I�p�HZN�Qn� F�G'��_��G�˻�f�s�ii�VV�>�&���Vx0���hN`y?�3��}��׀����W��$˞�ٽ)�~�3^��3jVxȮ�d��?�Ψ]�+T�g�*���9��n��;?�őpxҘ��T�W�cJ*,���� ��FC�T�F�=_��:9�:����bҖ8�Ô����t��ŪNu@f���hg����F���JO:GNTX�p���~�v �V_zQD鴢]EL�� &%���"����~�e�~R��`gY�|F�MrB�f��̱X�4U��-|W��$��m6҃�\^�>;
�h��F]Շ�Q��?q�I��OyPY@-dȟ�C���5H�@�� ����o�a�Q�R`��s���֖ρ�pwά���Q�,�ֆ������d��]��D�-5�pr��g}�����DhU��r9���YU��}7x�CXT��>�4����:�[��D�Ij� ��_v�-1�v��az��6���M)i�� �i�#=��d���9G8"��"�^�������!oHw�a�0<n�ӃT>�����y2��ML�|uKOatcr��h�}�(91�=y(��V�sD��R��YҢ�[8��T>����?4�6��&�AH�=����`>y���*�m�ݚ�s�_�&|��&cV���[�ǽ�Τev#�P�V�6�OOnK^#�`��-O�s�p��_�P�z��}5`�*�`��Kr��Xq��M&h|7A�W��B+ߞ��e��� �2=�<	�&���p�\���>�����������o���]�[1���{q�[k(mqwa̹5� �(��v���hrcw���ma#��⭝f�h��0s*D�/8�{{��f��MU�W�C��`�Br�Ӆ�~�D���'�I���$\�M��&�ݐ�R�n�1�e����,K̸��i8|Y��S�����T����E��c@�n@���8	f����L$)��e?�8���lH(|��d����
7E���8b��=�՜Vp<�4�+_�@�s5?�Wnp�AP���9�Nf�}J��O|KO&�b�h�W��K v��w�C�
蹭_��3Ծ�d\%���S/I�PL�2�0ψ�w7�z{��N�c]~�[�))���s�<ئER.�����P_ȼ>�v'd�V"_�F
���MZ&*k��C��e��Bxŭl����LD���8w�s�A��aܷT#���R�ş,ڨ��X]05��{��EED��b�l�VP4��F�S��6���.� �wb��H����H;�S�L�A�M�આ��PA��԰H�Ӷn_c/O3�~jW�a^T����.~��db�ڌ�^�\��`-�9��9׵��\��h�y^�?�\(��H �J�����g ��h��8����gǿdk���4�/<_�kƲl��Iܕ�����׽��u�,+дF�����Gڋ�];��}��n�h�K*8j�n	��l]���P��,��WMk�V��M��t�p�VСGQ�MӡDMN�����l{z���h$�W}C�y;n1V��L��1��ZV0���~�fN*��Io����5����9���W�x-L&c<�8�Y�g��qe\ԇ!Q�_��hJ2Wr/&�D��Î���݃sV� �� ����H�3�2���"cPv&4_5AK�ab������,A�A4�B�3=7p�@�)���6O�w��#u\�р������,*b_�X�ρ"uM�V�|O9�Z(��Q۹�4�4�=�.Lx2*D����UQ��	���$�E0�,�+#ɽGq�<����0A��Vƴ���:�S��w�ƈF�`"�	�0��E�b��r��t��ޅ&Wr�Z&��N���|��q� ����+z1pnpV?=����V����*�(�S���U"�����Z����P���*�7Z��l��3�ÎZ��y}�f��f,GD�Wv�������P;*���~��)�֠2�zt���LE9�W� o�1��h�[��Y���f��D@� �M� %�ġ{y�M�-tN�F@c'�l�^E�n�x��3&���B�j���JV����N�%�P�8��|]HgP7���zFb�6qhl�D�~s���С;{)�y��1 Ҝ�1�㗍)���H���e;����uj�����e�D,;�������j5��"�JW���g���s�C���Z�o�n���>hwvW��5 �jC�*�^��~N�/vї7s��[�eZu�f�[�����2�?� ��J�@��%��%���bj�r��q�T�r�}��&V|��]�9y�s$�.�B "�4���<���!σ����,aOA�#��ze1T�����I� !E�����-���Z�)�;b;H^p�kڥ��p%2۴�o:����s�4�����k���d�� 4�Y�Amt��&#ʻ^���YN��&�����i�x��B.!�̹��ŷ�3_�n+����i�w�p��5#�S���@�E��z�(�]'�]1�;�V�ٙyq#�o��2�5䂥0�e�7���� �d�'��,�j�`��'�-� �
������wu�g��G�U󿬤����������Xy#Y���<�%��SZ���àP@>��8+Nl�����&b �����N��x�͝ǎڮU�TX���z�'����i��\y0I�Zf[����}�����}��U��^�z5;f�K�(g����͸1�)XI|x��]��^P1&`� �.�o4��_C��,�^S���Kğ�=�(�ȓ�7x�<�Ȟs'5�ȩ�|`��u��C�Ru)�I�_��^R2.|����&�*�S�h�;�VĤi���"~K���Kc]��<�(YL�{������}	?Q���M���kQI�pԆ�s�N��h�r���O/��˛��#9��B8ڕ�qhx:pW]	�����n�5>p rm?��g4亍�{j��8��يqj����!O��t�nV����k8��a�s/b��F���2�E�X��G	k<���T� �#.�����Z�=T'Y�&���ݟ���6쏴A�Y;���Ƹ��u>$�c?�$��6��R�RY����?�I-ۧ�[N4Ò|�#LQl��@B��w�ę�ٖ��abg�(���J�@��Ov(��W�8%M�:��Lh��M�^��ox�}r�� �{yF_�Ҙ	�>��vR�����R�B�~�.0�}$��O��-K����VH��9�����a��� �l���&�� ��`�ǭ ~a���Ṭ�"����$H�)��վo�lFaa:�`0�Wȃ��1=O�e�4;p(V^�N��\�S�G�U%M��0;�B��<��B�v����Ź)��ԏ���&<#oy�������F
�~�֍��hG�c3�I��!@o�V@8����P��YCF�c8��k�כ�l2���z��{0�\�G�7`W@D�s0L!�]Xu�`���".62K>!�����M�3�d�To�Ӧ<ES���ʘI��v�����*��`ǰ�'��Q3Bf��q.xY#b�6`?�ǥV��T���?;�B����P���}(��L��5���߼X"e��ʁ�j����G�z7�S`%:\~�>1B�X�=aJ�e��4!��ZX!�Ơ��5o��\��B14��3�&�3?��"�� ��t1� ����31�L���U��t�ZI�a�;�`(b�ig� �Si	��.vX��1cʤ�9bF`l� *�a�k.�Wg��kʾ�QO�K��i��w�џ���`	���^����S�O�x5�pd�|�"'�q����#Mu�����C�L��K���K�\n���0y{tΠܥ,��6C[�E�?��E����M�8hlTD�G��]��7����e�lsv�\�h�~�[`"�iXf	$4��J����7�pڥ��`s�Eh��G��������hZ(7���кa�\��ɡE��@�8���|�T�����D�89Լ���!{h���:$�`���"��:�O��C�^��%�c�IJyq�ckT<� �\L~�d��aw2����T�i��=U�I�X�ZB�â���O�lP�'��N��ľ˵�m��!2�p��MTY������)	��&iН?�k~�q����{I_�TO�ý��SOG�J��P#ʐ�9.R����<���-!^���Z$*��&�MLb8�'Vo�M�fʢ0jZ6�+��`����O����_�� o�W�m�H�_8C(m��{��FU�A+b�Չ,_	�K�Z���f��:��^��@����9�s�%c�0yTX�\��id�y�sO���9'.X7�~]a���q���!�1�e���0km���r������q��X��#F03Gb㗮�9s�	��w�e{V��,����f�j��--WF]S������TFbǚEѝaw��:7~i0�x�_��G�!"��E�_v�YK��{+4�����=X$�6mWh�@�?��l]�7=`VnFq��k"g+��<�GW	�PFx ��L?ɺ����������!�4X�I�hɂ��T��+��U�vMd��&�7<�8������{�7�y�>�~���P{���e%��:{9w��h]f�n�1j�P���U�����\�1���bZe��t��
�?��/-)���e:{@�֨-�>]9A���[Bhʝ�+��4Cs�m̷g�w�ɋq�^{�B��^���#��#g�u,m�za����o�⩟F�f�[b�"���?T�W��W;��L}�/z��<��M,�'J���$�dTD�4�ocSݲ�`go�I$}K����)�e�(EH�����`|it1Q,��9N>�r1�Ԇv��ep-� k�ۏ�g�m�WZ��b����r�ș#������iE���E_�Ƌ�����o< N��DIkU�Akc�R�%�������κ�>��z(�����ͺn,�`	,�'��*�1%�hq��I��A4�Ձ�	�$�`=M�7��w8z���y��0��X�[�ë��;��y�@΍V�HM)�g~�_/����%�ǝo��[D����T��������z��F2����#�c���i⡝���%J9��<=H��ŉ�٭ni��0P 5{I1.>����G���R��y�R�nx�?�c6'��R�"2=�hM+D�`�5X^�t�'���)�DE��#>���͸�V�eס���?ͬ��2Ζri��;}�&{n"���m @,��XK����}ſ�G���o;A�x����������På�)J�qXH�@�x���^�9A��p�˯F%܏�:�Xm�.���D'!}|^�����2�Ր�_e)n�p���<�}\�:MLFJA/=-l�M��k���P!R���`�j p�s
$��9�D��&a������Yxy���LG��
^فZ��\�Y�ߋ��rTK�k�l�X�=<����c��W�XD���'�8�ڣC���1��<
K��F���4��&�f^m�3����_x!:[�����������Y�6mη'z���@��ى��Z�p���DP喔}�Y>ąˁ����� f�*4?:�n�[�=��@j*��Z��DK�,RXP����+���J�V@�4���CNe�@�5o��n�c2��n��U�A%�P��tk�³X��67.�л�dY+Zb{&�pf��^�'a���f�g�}f�K�sU�-th ��W�O���xp.-$=�ͽn�i��4 Z*?"I���o��ԁ���ϖ�Vfh�����"�NK��w:8ܲ��} b�.�g��(	�=+��n{;��ݝ<x��L ?�f����<_caa/6�h&��w����w�g�Z�ʢ���Zkn�7� �d��1�jA�F@�#eZ���o�Z)'�0�#9KH��T��o.reA���\e�s�%m��M3��_�=��a��W<>���g�D������� ��}��1��p��ͣ ���L�u�X�y3���ԬZ�s�4^p�Ԇp��&��1��_
���Ux�8If/�^6 Fl�Q�"�J��S���N�?o�S`���`&��rFژTSYӧ0_7���F`�:&�y�r=��+H����Z��U���
r�H�("���K! o��OU�#��Z�j�#�*sF�U7*�K��3��~cZm��d�����U8��5�H��6��߷��{�������P�9�%D-�[TF��Y��2�`�(�N��� U���Z/��%����Ŀ�7� ��W�r�d��G,O�*�Ҕ`v	|N��ET�VĤ?��Q�ۑ&�h�`㈌�u��?�n��g�����h�70����T��ϑC��c��X��IH���L���h���mі�+�dAHGX`��,�^�8>�.H�G g#̲�Z�t�y}���D�(:�	Wt�s �/.�ߚ�K�������({�;�f��>"K.;�PĖ��С�n�׋�^�kF_l��;��+��~-S�b'+�I|af�L��`ye3�Wȃ㫿84 �DD*䣴��*<����W)'^���@|�ع:�t.�C�b����������wQ.��=�������@�v�?U�Z�{}8vsA����ONf&m`H�cMA�d��ψ�_K�B������*t+�� V��k�Z+b.t�M�0��U{j��l��eߦ��-�-o���jcW}�V�Q[�y�)�=x�:��+��F�\m���ָ���N�2�|r����+f��\��f�K�Ұ�w���K�*�@�'P���}��㖃k�} ���Y�h�O[I���Mq��.�ʦ*V��EU�g�qW�Jw9���:f�~l^ُL_�SvXl��{W�Ɲ�����Nd*���rk�t8�]+�N���yR>�Wn��ƿRn���,�H�v�Vmre6_�T�B�65�6��^�d��s0��z;$�g_m:6dK�Y�v8�)�-l+eܟ�\����Y����쬲�ٞ��v⣫���~��+��	�l2����W��K�fG��Dn2l���iBspa��+ev��_�?*�J���P�p0�XR����&�$�g���);l�v���� )���GH9�h�ݾo2��?�@*���6��G����:%K�����Ʀ0J�N�,O-�sM7^�+/v8l��C��M��%~�]M9��E��RI�CI������ߵZ�T���	Yډ�_���{��q�6����5���o����A/[�'�Ks�ƃ$� %��)#��2�I��;�dgBB@f�����$ :�风���<���t�����u�9�h�}�Ѻ�i�sx=��;}�o�J���&­���pXY��Zݥ������7���-�- ��_��� �r��'t�-�����3�G����:puw��H��HOL��g��uV�괿�"�LT�qR=�fW���I�����T��J���S�w��5�{�[q�vxy���������g*�DEc�nQ�wǵ��^��\�G�l�2RT�\�j%�~�u�7@&?�*n�s$[��y~�x1�+Ɲ��eAl��9���,�H��
8C��lS5`z�rɬ������)��h*d�ƽt*�K����G9#y�~-�t}S=�?�`���P��Ě|L'����άQ�F=�O�Pӭq3Z���E[XH��@#D�F�u�A�,l�[�������.L�V �o�|Nة_�*���s�:�¡���/]cTǣ�E�Wy-�c�
���Aضc��_f��;�_���]��>�W��|���7,(���F*���]��H���l��l����f�>y�|��|�)���Lc�̇ޒl��������8[�\�p�������ٽ�C:�]`�I���G7�l�!g�.P/����%'|U�&�=�b_Sl��y����='W���8��2�G���+��'��la$��$�(@B��0@����AY1;���vaVf�oo]i�2������wƜ: 6G�aaT�u(�,1,y�~�z�:�D~�&&�A���Qv�Y
p�
F�tOب����A��ْVb
a��f�;R��d��`�y���ݍq��h���g����<��Fu�:Ȋ-yM-��bU�όc%Ty���ja�q�_�#-����pG?�iXd.�3��5���}00�GaO��2��/�h?�e�_A4�nV�z�:}@�G*[X�IL�F�â��~c���ղ�%���'ڲA��q_���G� L	Κ��dP�8�����7h>�2��:i��1!��d�S|u��T5@�^�������)��C��v�b 
' �޽���AT���6ҝ�M��Ѽ�<�qY�4�]/lR�9!�p��e]}`���x�{@�y�"q�yy��(�{c_R:fPC��	�#!����P[�dc�ـ���ՐX�&����ݛ}�ʧi�Uk $�쒈=�t�X��S�FHb��|����:ئD�4�C��*D��^��2y-hM�)��Ćq�ю�y$Yxrm�(�k��J��R%�������<hL�D 7auH����Ed|��8�͓�g�����x����G�s�X���@3kxP����D������"��ɠ��~:��8
��A�΢���]��E,.�)Ca�oY�M���7.aO{����ۏ�5i����rA9p�$��7�[�f��sb;�57f��k4	w��Z��r�(�d�g��-=���W�B�K6���Z*�f�.˕�!ǐ_.�n�JSQ�awV�	��H��k�n������PQ��I��U�q��������k��!�$��	pL�mCl�]�*oM�Ben��N!�������Uw���	�����p�w���Z��Cc�կ�o�#���믥�"�m���.Qizڳ���j���"��]�wM3�[*���@��pP.ew�3[[��hG!�@j87)n�G[2(?o�^�� ����yǷ�lTjm|~l0�fP|��p�>V1�uϚ�XQy0�����Q:���,�T�DDS�O����nś���Ë����F�g��C�T��^<�;�Q��Q%�|������?���A��+C�8$�q:v��:f|���)��B6*�w�S|��Sw�=)����#�)B���J	Y�D-���~&�$��Yp:����wO��Ny\�A���,�Z���v��vN�'n�"
px2m%���|�?����'�|D�>n�#&��q��8]�njx+���'�d"W ��G��A�? �˨Yc���a[�	�Hn��y/wF4�+kl�7��@6��O<����0��}Zp���a:ʚrB;ܳ�O���|�E�t G`��$��M�eJ�FU4�î{y���F�v��m��*�xb�ab�*a0_��r�Wiy&]˻i���l݄�x��9I�y��v��Ai�k%�hxa���٩�O����yi�9	|Db��h��i�.��`
 r��Q4���p�>Ml*;$	q�����j�Է�ni��tD#�sh�S�y*Yk��E�����ܰ��_9U�3����+`�t{B�@s6w��[�	\.��]����)�j-u���u������Q�݅��|�l�T�ͯ��⑽T&�=��1����ذY�QFuKǿX)��>\0�����M�}LK)ɇ��U�A����@��ux�o�,���}�D'�<�j#Q�n˔�G�G�d6Pe�GDq�f��P�=�?����e���k���ՅW�&5� ���XM�|A��Q�@���]�ACs�appվ��#�i+^˞j����]9JZ=ѱ��S!�J 3ۇ)�<���* ������>��rl7���������F_9�s��{=J�a���u�z���!���+�6�l�E�4��L�:��-&W��6�l��`���w�&�a���jo�	b7$�ܠ�5�v+)�	�h�U�?e�f�at��fa}��jÑ	e�;6C�p����K򿷳f�ŨG���>;�u�L�n5�ʄ9˺�rA+�G��4)�on�~.O�h`���"J�\q�N�/��m�T�ۀ
	K�z�N��X��Z�@;���[����s��^ k�g\���'Z��m�/{ĕ/?������r�%C�!����P�G,X�/���q<�ħ�N�m1A7�{��Bf�xV��J���+�����J���J#;�cr�=2���QD/F�q$��F�g^
�6�d��<��n�����?��,Ņ=ki���+�G��umo.|�rG����65���豘�ԍ)o������+�P������`㌁����[�p���}�>���ī����'݌2x�,��-a]<�%l�eko��D�Y���t'�B$ì�_���C�\���(�=H���3 {6$����:�6Yw�g�8d_b_�q�7���Q���*]�.	�$��^p./0z[焖�:�(��-�VJ���7�C��J`RYT�M�AeI���^��Rz�^���[= �4�ֲc�&����%h��eB��k�9nc����,P��Es
�yBNFk�Ձ��c�q�GYt	H��q����a�	>B�%>�Ӊ�,��Ih����A�̻�=7&v�$��-C>t��}��`&���׈��jy<Ie�@�[���h��($�B"#	[eh,v��Y	�K�L�@'9Ld�~s��d�jnvVu�Z�B/��¡������:#�0�d.���p�~���w\�4�uzR��*��|�G�>K����W-l򹠂t`<�5��"����_pZT�p�~���oa6VM��upF���p��lp&�v�C%��Z�0�>%��?�j<;��&O/��L�;��r�Z��8�Q�Xč:VK}�_���vu5� !7�z����U��تjdl}и�� :������6�?�4���-z���ɑ\���4_�%w7�{�r���{�^�����mmH��/H�ҷ�R�*���M %*��lA��i~�R��=��Iu�A���L��6}q|3�S�ݾ[�śy���# NB����B������V�uّ�;�cL�Uj{MaL��t���y�,XW j��n7��C�&�%)����E)#��U�/���n��(��v����Y�_0@�0��[b��[�r���_�����5�x�}�9/+K�A}p]���!�Cԓ���;�_QԄ�o��&1�i��r�A� �ds���팈8���D�9�N�����<ߒ6�9�V8����</��a2��7	�w��8�8����t��`������jU��b.��#�*�Lf��
����
�D�<�N�|�f��tbP�����|k�7�5ju�6yA�F=떥|��\z梑3�x�L[��Nf����O&l�#>4 �����UJ�-6���-��[�K����8��~�Ѯ+���?���~�|�Nج�ctC#�
���Я���������n]wD�[�z�G��m��t���2a���t_t푘���&�Dg@>�b{�����,��l=�D�8�Q-R� ¯O��[9���٦����vȹ�����JF��eѾ�21�e�^ D�څ^�E���%�Y��ސ9�n��䠛�\��ר��vX|�n&l�c�І��ŘǶ�,��B
���������:&QzCh���־s�Aϵ�hy��.�U��������CI`�2m�'\�AKD�����I�|ג�@6L�h��dO���#Y����QD�:�����2�fx���%� ̀���L����k��|5�?4@7L��ncN�8��g�Q'@$cu�{V�?m�@]twr=����X�{���n&�!�[�o�ͨ9�4� �r:��C<.c��i�K���&��`U��$�>hI�7���T�Q5�"��p{Y$&����vx�f�������`0x�g��5�wH8d���jY8��眾��DD����X�apX�m�S�$�^"52l�f�nZ�G"�T�e���F�� �����z,� `6�W}�6 ��s+ZC�9#1��d�J��B�}�<�Z����ٻn��̹��nt�.:�w(�/�ޔ�(��緓��#<�i�)���kR��z��5��T������g���(g`/)E���;���*�L��$��`V�&��wcz5ج���69��b|iȞ���(�Ci�j+�|У�d�\UW.�� ���k�q�>H4`9��{�dr��6.�\�rb�R�r��HĔk��(�cK&�+�.�H�<\�ڪЎ����D�/�N�~k�I���� �4�{$�=�6��\�|�"O�kS.]�U4�qY�X�hX8�o:k�or�6������Y�k^�8��ۛqq<7r�Q�T ��h���}��dݻ��IK�2:��K:�%�i5<�3�r�	9��v��"��C'�
�2-��%Tt�\B=V
M�=�#m�L5R3,5z��&R���F�X;�F�:���f�o�θ�h
~/�Z�;�:"�M&��K�������<�Lʯ�+k�_�	�dC�,|���|�������'��}D	���OUl*Ò^5-v�H��B{��h����H�_q2 J��j ��{L'�s{G�W���L,ÏZЩ��z����a�����q�u<� �	Ք�_0A2Ƥ��[T�=�	�lw�c��63N1P�32Y�P����$}�����LD�\���@��ciVN���EZW�;4'�+[�`�����6KY��1��-A[�ޱVpd�gg%�*2^�t#Sd�Z>*�UԾnK��R��Q�ܫ������1L8�^��(ʒ]��� �ѡ^j�E�~Ι1���w���uh�sa���|~4��v�r���N�g6���p��"n
�L��ԑP��21�n��1t�@�/3k㭠=*��6���I�!�e�`�()y[��v7�\�q�3�~��%禸.����� C���ħr��~���r��g0�ˈ�B gI��5�5�w�� wٰ�fp���M�#��>-ZF�3�]�Y-F�oW~ߨo�l��
�H�@S�d��Ҫ1��K�W&��$�7f�<��eR���Ni�L�qL}9Ϙ>�I��I3��]��\�J��G���n÷���j�
�ʍ�PX���Z�f��ɧz����Z��7��⏀ٷz�4���7�U�S���ݏ�� R�!^n���!z��s�i��B�rk!I�n}�o���m����G�x��tb��|4z�y+�L�$�|�z�r#�ޣ9����Ӎ:�a�	����C�M�,T�K�w6��1�<�����ؿ16�z&���/��k��6����}����G��7R� �I��g�J�jL�� '��q�s���PNOu��0�=��(Iٝ=�P��-�d�M��nd�%��g��W�K���)�9�w��^�����;,X����8yO�X�1͇�a������f�;�,�H�q�U�9cݓ�/�ԓx���Ւf��]�^�`o� ���c���S�Ǘ5G�<7��:��6�*��5�u�ί3P�" #$'��<E/�=5��rcg�J�=�"Q�2��>���-'�R�CiY�vL�Cz㑙#���>�|��QY0=�ߥ��0B�C��Q�KAJ��v�0mO1I��W���=��F��.�>�N�F��ҕ���A�� L�@�2�
\
�_���t,1�>��RnZJ���P�W�.?%O-�,,�jm��K�������P�Ǭ#J��hnᢅm����{�6X�|@!u�Ň,��I?��V�VI��o
��C=^���X��G��������8~��@cx<p��̤�k�y�4�����D���;�N�PvA@���j����:h����溒${R��rg3u[X�ᓥ�C�ƽ����\\�uXv$��v�;<=l��+ZW����]�~a�n�C�A^�rkY�u� ]=ES��$3�O�4_�U����ޘ���\����S�z�w1����b������Y��ѩr�����ܵ^�*M+��|�+vȭ�m�G�k��t2o��sL��ox���i��4&�T{m	��XOμ³V���䥎�l��"j��`];>�p
.�/�D�*F�H��s��%f��J�g�=q%�ʼ�K_�8ֈV&G�5`����{��?�9޿�UCy/��-w�l^B�e|.�3�P���c�b��_X�M)/x��	�s��+�9�{+Tn�p�_?Ů�\iY̻�?*��-��9q&l��*z�?�|$��n<�^�]����q�X9wPUZJMI0��#��C zhنCn;!%�n��?^�V+<Y �9j6�'
�)g�-��2_�k4
¤�T�*R� �eW(e󸊪\>�J\$tT��� N���������F���|��.-��S=�J���>e
OP�+.�ٮ��9���v}��M���t.�쇯�2�0��\� }��Zhp*� ��C�%
���&ݻ��k@��
��">i0<C)I'?��a�XE�F�L��(!Vk'���#8�F6vfh��ϻ�p5͕'P/�X�Q�jU�	j���^Iv��]�8��J�.�o�Ҹ��M�"��x]X�+�4���j^��9����k���-j��4�i#(�Ͽ*�
@D8�VZ�h�G��GK<��<gՍ;F�.��(��|��Ĥ���`����YN�FT�
-|i�yȆF�@p�Q�&Z�B]��t16�V����$P�q��W%���E��&�����T̬�pY�gL�^��?dèn�E��L=Jʝ׃�!��C����Z%����X�3�yh�62>}!��j����"��\9�5�/?�w9Y�s:8�}1+zӋ%X��ˣ_�c**;�Yy�4���I����DiMM������7�id����G��at�յv���F�ֲŴ(�.�d�)z�9��3l���>��o̰_�Ѿ��q���:q=MٌED@�d�[�8�\��w�7j��T�m>x�v4j9,y��s���� ���.�Rw!��8���p�BDzf�HI�څ�wW6�B���t#�v����S���)5�7�ȭ�|���>y&��ߞO�4�>a�E5�?���m�<��zj/���"�y�Hr�Ӣ�����y��7yt-uO?B��Zʄ	55��:��$c`l
v���	���p�4��gou�U���jm6"ϕ��I�0���G���H���)��ʃ"�x���ы���v]��z���[��Ճ���JՈ�#G�"���k�i�/s��*����.�W�w_����6^mk�����{��I:c��8pd$�/����=��)q:7i��H���E0���
HZ�9�<H��7�@j~]�`'������J)�~+irm�I��|��!C{a�"�e/=$�$ 8���9�S�L�2��!�Y�ɖLnol�>z���X� �@�>�6x�z�����;��^m�� �owz�6J�W����6l��ҝ����]����KqДrȞ$��b�-|�	�n�ܦֶ�
��	.��B<�KHbM�d�ܨ��d��PL��K��|�%����Dx�'ݖa�Jٛ?'4?�Q3�蕠��T��L-�A7f5�x@��s�Db{���$�亄�U}�k��+zH_�w�}��m˫E�鿢�(1z�{^T�%��g4�B��Ay������?�.���p��9��dЄ� /���>�h�BcR����ISzT����
<w���Τ֚+
�'9.�-���ԕ"ZO+�M�*��ݯ���`OR��G��S������J�J��Z���	s�N��Q�{��s˖K�����b�_56� 	�����N����̂x:Z/�ErȠ�g��S���~t�<,���^�x?��p��=���V�J�&�4A�M\L�سX"��3��p,�[H��4�37x8�,�,l�w���IgV��3��v`�:����y���4"Z&/y�j��ڃ�����;i�I��+�DZ��8'�-�6���&v"G�8wI#��>�yP�g#NGYt6����W؛��=k�ŋ�@��U���R�mx4\2Iwc-�U��:�uX��ߝ�š�3M-?�@������Y���� X� #,�7ώ�2�e�_ᤂ�X����*�@�"��˖c�����oZz����".P!ݶ��� ���26h�!��m?�<|�gj�		��5�n��5@���O6�w7 D�~���V�j����d�'�E*8 �5�*4��T@ѤT��}c�M`	�Gs���f��-�3s��������a� �>~B�����z���TC�)��:�Es�7]dc_�v����)F�O@
Ǟ�D^��l�JJ�U�_֋,G$�[�p�k���x� l���U*Ѫ��}"��y���Z_��v��WZ�,�ēt�`��mX��`I�-9���T$9ﻑ�@�\C;v˜H,��y�}���	����j�Ӌ���+�FN�N/:f�VU���EIP��o�a���($%��v(9u:�{@��f��D�\4��Ԯ��O,0S��vF9tj$�6�S	]����H��Q������"*{���V� ��-L')��ܼ�u
��pͲ�w}��GlRvqU���v�*�J�H�?t���m2�ǡ3�^�8��x^�C��l���3��El��QI��v26B;J��f�+6�L����b��+9CA���V}ŝA�Lu�FDm���~]���p�H�#J��
Z����gƓ�CP�T-8X��,��T;�Q���;��
jz6�E^�V�."Pe2O����Ã�BR�z��{}��k��4�\O*�mz��_�3*?�	�>�8�Cnal�G����`�Z�%5U�m�JG������W�ۯPl־#"l����%��)Dw��k���+ 4N?vݵ�Z�Tj�@�+&I��.�s�k�J���v�P"B&�`�*y���|%1,Ajn�E��6�m�P�
����8��";���gf3v��O(��
L�B�6R�u��{�*��fc�q��KM�H�+��ku�|E=�-���&
�-k�_H��r��C3�:�/(�e�=q��^�0����tu�h;~��4<#����$����c��7�Ή�h�[��g��Y�H���R;�!��#'$���~����P�_�dz�g�u�C �lk�g�J�5R�p��R?8ZW+'�N̔5��m>j�F=��R�DdTr� y`�"5^�R����p���$�����"pu�Ǎ��f���[e��Q-!�a|ܲ�	�>��7U6M�Ju�>���M�O�nLWI��)4J�E�귬TwU_�� ��@މ�!�I� ��P�Q2|3�E, ��Fm%���0 ��Ǩz9�v���!���ʭ���Q�6���	T���$4��Q%-<�ā�(ZQ�=�2fAy�jvGM�����/!�(�_�&�y��a&�33�/.ybZ�n���M�|!�n�6�yP�N��ꘄHA�FE��Ί��D�?�8��\��Rt_<��ѧ^@_m�h��by[f�{:����i�೐�b��u�*�1��JX�H���`��y����*_>)��*n>�GĜ�������^�N䜌�7�6���1]�8wEX(qJ_�����6�d�^@��l��e���XQ��.$1����"�dP��~Է'��rh�TxNB��ȹ����Q���;r����;���ip�n�H�GB>Z��8���·d!ioò7�����}d+�,�2���*Q���+&pu[���2�q�����?����no�e�&��ԅ*<0��y߄D!f���N�����f(ӥ�1�����`�M��
����M�O\x�kX�]#��6�@y��د0�k��ԏ�+�r�4I�C^��027�3�H9�Ԇjut�s��	gXK��e��G���y�2�E�he�	{�N�<i?��rc|�]2�����H��D �i}(٤�P�~�Rq]
���\ӧ�v��e�}=m>
q`L�A׫���#�v��-�8��UX�J�R�ʉ��[[�|�7�G@�ʵ���d��y��tU\�G���6�:��d��c�\�цh<�u��H����`%ɖM|��+�뒪i!�%dJ?��Ɲ�G�ZJ��^~H:��7�vw+�뫂.��:��1�,H��$]�������5� ��x��S�f2j��{��x�=�8c��� ���� >r%W�߯���8�+�=@7s?I�sL�)�*�sG��YӾT��_K��I���Ji���xcu�20||}��nŲL�
};.xxyu�/Az�l󤣮���kͰi �##*�9��'c�^���ŗt��Ӱ�����w��*s�����)H��;�۞��,$r-�֖(���Ͽ��>��w�s�����6�AU�����y���=���`(�2��m␽���Aﳷ2��`zh��u��O|��C#$�!��Kv;p� x�l�
P��G�vmH|��jX���`�+8�ޝ��=++�*.�|N~99�{i��T5��v�@`����ߎT��0]�j2ڍ�
S��?�3Op��?��;kN�z�n�4L�ٞ�=k����I�d��d�V~�/�\��+��j��SQ���aDBSs��fc%)Q����ZUiB�"���"���k��@�uX`��ZI+��0
>����|s(�hh�g4�%��'>+�i��b�o�P��.�e�Zq��G-W�\��<��p_�"`V��������CCp�fh����)�k2�nGWk��6�����e�?s��TW�3�ţC����Py5����������;-#;��{�v��f�������}���QE�Oa���'le�W��\�,�r��t�)r�:���yu�@��>��4�v4��g��[��8K�ɾ��
f�"�r�4��6��wJV�?��a��B���;��ry";�!��d6���/�L�έ��
 �j�0x~��:�b�0�D���v����Z&o;Br�7�YO�{ը*V&�Оwn�Ґ���Wfo�ڥ�'S�4�K����#��|A��[��'*�I��ե�t��+CK8�����H��]�N��Y�;@�=��cv���d���y�T���g�@�gK��rfW0q�Eh�5M^~ѝ�g�;5h,��\�	
�V�^��= N���k����s���
�s�	f�V�V~���mO�K�h-q����**&���S�|0�A�6�D�����#���܅��E(rڼ����$LE�ԭ�"�yp��?�MD�a�;�wL"�6���h��E;C]�{��z�j�e)"�����2)S�Z3��V�Dp-;<��}�r��(��`i���?@̚�,��g���oV߀��S/%�ѓ��.���+}m�b�#B�X�8��`���}"T�6�pe/.�,��<;z"A������j+q��A.�n��~�φ�줦�N85��,[8��v�E*S�|o	e�ʤ�Ej�N�8��=���!�ӹ�:�qdh�}ZN�ز�������u��r~��*�&}ŗ�r(F�4���)o8*P��7,�Eŕ˭��W63w\+�jB�pӒG��V�KwWYEr�G|���m���P��m�\�&�'��W0F,���73�đ��t��m�$�ݻh�9J�_!ţ* /���������.�-�:��}��0�v-�CUޖ�����C�o�(E-��2�бfeA���i�tɊLBmc�����6�
��@�?��&�ĝ��ߋh��T�g;<�����c~���A��s�4���ї[l�Tqo�,fqs�F�B@x��M9�[�Z� �����@���r>���p3S����Fj���PCg�׸m!��.��bL��0�$XO�,��p�^X �f�J���P6��&&��XZW�iw�W��U#�u�e�aص�&fQ������-ŉŭ0G�Egwwd�Xa����}���C���^�������H��&d�-�����.5��!�<\ ��.DM���2�I��C�.��J��!wJ��m�4�X���D(�D.UV�?�n��3��)�ϓ�8��f�27�u[2���@��V��yv�?v	��r,6��ݸ㤘r�J��ZW��Cp}J�ξO`���g�֮�ޠ�� ��~���Z�Y����Ymш?��j�X��X�$�6���n$�4(��C��'Hz���R�s�1:�����gWnHx9 ߓ���i�
�[q���F�9�_ȣm{0$�-f�`�`���J��^"��c��O���<<��纘͘Zsrg[UMX�+n�A��П�╝�fQ��n}�
ON#0Z7%��SwF�����_Ķr��V��E $�"�:ѱ	���+7*��~�ݭ�^b3��-_C�rDy���.��aXl43e�p��;?�@�
H���V� j�91��g���{�^e�a��ai�꒛Ex���f�js�����(#n1q�%Vo����-�����(�(�L�����>�Ӊ�!�іn�'fK8/隉�o���-��%޴b`�H�g�8%^��<��<�:��&��ɋ���v����$��bW>b��/o ��(��\�@ݶ����)��������>Vr������_��Z�T0�PV���e��՗%�	�:�7����Zύ�pW���� �gm�b�W�;C����"��)�ޡ�i��x,�� �)訲�I8��A:� �k]wW7-x;S���<��1��Rxr ��EJ'���@4�-jA�q�o9����$p�-)��`�>��
O4��nГ��WUu�����������q,7�$/�B����N�����1���`���D�.�Or����X� �ߊ�!x4gn�2�y��NF�3�l��2,�[:����f�ײ�Ιw�B�X�O�<}B���#캼w�����w��^V������_��O��z5��3��J���ع�LS�"��f�g[ ��,1p������V�?��gI�2��1	�R.��=�V���F���H�ej�IE��;Z���!�'R�M?a��@Mf�/˷�K1q����ٽ��A�)q�]~7��{h�X�3��Ir��2���h�����nF�	5��O뇳%��c�6�)�����6@��Px�W�5f�</Ժ2�I��U:��X�W$ ;�?e~�\�Lt0e�_F|HOe�Yl�_K�{ӍŞo�5�G�~�7AM���D�Bp>"3<'���D�X���]�ȆB$Y�!-���^�4�1���$,d���?=K8*'�҃^C�ق6R�܊a�J5M,cs�p{�F���y����|5�b�<�}���p#´�v�q�b2��`�������~�G�;
[��s��4�J��r�I���j1�C��n���IQ���e��'x��N�-VsP9Qg����mV�1��j6|a��v�ùWt�]*R��V�~�󣲖����
0�/k�)�I�P�~Y��ɏ���c�5�Ű�K��i*W�Z��O��4��6�6����"(>�%w�d��+�8L�H�U�pB����뻪l.)C?)Ri�$��!��7�����[��K((C�E����3�kj�����o��F�J����ݝ�T����X�9jk�|@�?'�|&����!��ݒꝳo�2��V��O�/BY<Ш��)�$��(7G�^�����sM�ZC3��=<Q���,�o����Z)�ԯ��8�t�t��_�y��^*�T�'VL.�Zyz���0Z����2�����'DV�ʀ1�k�:<���X"}�5	�@�!����z���r�E�Y���z���@�%�H�*�����A��q`N7�݇���u�}Fd=:0<�,¬hr �Ƶ��2F�d�����ra�*�+2;IK�f���=�KV˫���p��݁�A����u�K�@���c�e�N��t�8�G@pa���5��i$�F��.��v� ���^��)�����w�Ӫ���"yB��	<����C� � ��!k�5lj��8 ��0�U���Qm�Al�ˍ~���T��u��m�)��K�+��)K<J[X���V`���Ƚ	�SV�z�&"�-�Z�p�ّ9�F rJ�C�f�ڒ�kc��%'lS���ww�� E]���Z�`l5�W�]�_�,�M4��ჩcd�6�c�>�x�>�^�Q���Z��@ � 㭾�UC)ʡD�\@CP���=*���;�*?)
;&֓��M��C�B��L9s�Ĕ�>O1�U�
��`��p��Xg��V����%�P}w�Į�N���Id�Ř?
��i��W�3u8p�^�#��P1y��j}�DFCa�������^}/�A�i���`{Ǳ�X'���+�άΌ盛h���"�2�DHj�����e��o-�>dj�D�tmR�y\���b6Y��Xi�/%���XO�QVu��.H�Ϫ�;۫5�2�'�v?��޴��Ɋ�*f��K��8�#@Ћ@�JT^WJR�b޻����j7�L�d�O�F�;k���oM���h{��?��7,�;�!mE�Kj�)^�v!a�v�.���~�T�x�v��x��8\�\I���p-t�=H�iv��Kؔ�}0���,��р"�t/�2`aHE��$o��HN..{ʟ!8ãW+K ٓ_��񉟻w���0����\�����O}v��t{��������BS@gA}�^;���3�V��2�D�΁�̄�f@'���ڎVh�q,�Z���]V���v������J(MҴ�o��I���k����Vg��-��nR��z?��G7�iM��<D��״	!�3a�((��Qh���/d�*�fP�ʅ�ٷ�ӹ��U��L�ϴg�a�zP�|�+�}: 8��Vp�(=Q*�I5�� _�	��`K(*�Hr$�>M�I�v�+� H}
��@�:�$�%<���i@�O}�Ug�E+u�C�X[��R��"�o\��Şj!X��&�a��)?�ߥ��~�ک��]~���_葕n��Z�'��ƕ�ACBÊQ�r[��U٨�H�b�� �&���m^]i�����v�#I�P��.v�Kp<��a��6raXV���0΂_Ē2V�4�p`��VU)���:�,�bO�3g�g���M�j�a�3���B�R�S��Zr���4-�'d�J�	�M�tQ�6�u�tLKB汛��`�9t�����z,_�\?�u`2s��]q�nŔ�t�O�7Gڱ��mЍY_uh�&<�媻՘���򋫤�̭x"I 6G�����l1�\�U�h������� �A���Nr���Z]��3N��/S�1n3⋚"r��)�h?km�C$���ܺ����o"�^�H;�=Y&b[���i粦ic+5=�8ёo�6ݘ�|^�.3�J��/2���y����&���t�mȶ���˕�Z{��'F~`	���{�86��d�p_��j�u�'�5�
C����l �P���0��W;�*U]��J� �0���|�ZQ�@H+���?F�zl_�N/<HX�)#�x��Y�T�+"��<Y���9E�J�Ӗ�$�T�P�i��� ��Y�	h&�N�j���5��<�J����Es��1�H�%�Ag&���ҳC�/7��8�|5����@v�;f��1Reߟ|�tc)�Y
|"N�'{�岔'�lГ��`�V;؅K��l켉K�R.��T�����~��m�Ʊ3�n��Z�E�\R|.�v�� �ܨ�^�0��k1��K<�C�Ƽن���wa������������9S&�����%:���_���2�-����A�A󓻴]���p�4bPF1n��;��S��z�����X���`/9
jc��H�.b�&��巪:�� oi���'��p\��?P�P��
�5c`�ɽ��(���`�Os�{�`���H��)(�V�)�@ r��o���uL�I�t�墀0J0���x�Bn`g�aP��s-}�`�ϫ,����Y�"�S�,�U��ya���*�5��Z$�vT>�L�E
���WX�_����#������d�̜�n��c��A5�8�{�&�*{�6�q��
�m/(e�����g�ճ��$�>�f.��I(�I@�I����Z�$�?��4�æ@��|۵1)�j8F0:��/+P�S;?/��p��¨g0��R>g+`�̑�Å=�Ukr�{���&���	'"��v�ݽ��s�[^E�J(P��� �S��;2@�;j���8ግ0�"�3�ː��oVy�@
��ы��C�ld�F^i2Ғ�C[��s�o|��(Z��D��V��������{�$��í�'�9W�y�q�x��Q�/�S)�Oo��`�\)M�ۑ�n�)0���0�<;�ֲ��]XQ�����f�~�[~؄%�/`�����{�s���xP1{;D�}m����X�\U3�a:������섽��5��, 쪆U�7����㼜2L(6�� �pr���"�3�-1�����ͬT0���L!���=��Y��@Ia�Mv�j�[��"�� ��p��!�J��5�繱*���aRE�~mL���:�I�eX��E$�6hFcxun��sR8�4-��ȿ�ΰ�K�
z&�S~��2o�x'�خ��E(o/�t�����?��2�GF�S��Ax=k�|��$"�A��Y���{^8����z�6̿��+G[X��NV�h��a�ԁK���	���Qƾ>s$q���xQ��MZ��a�oD�&0��C�W�fԷ�/���M��(���S!��ݱ`�x��Xo�>��3�^Z�3D��*$)�-~$�6ؼ�o!���b}����1;�V=�H�='��I��氶�WJx�0Ό~l�����	����-�N������jy��:x}��h����E���B�?�\p�K1�=��3@�.��S~oE��piL������Ws�E=s�t|5ܦD�(H �";��0&��/B��`8��P �삿|`-#'2�����S.W.g>?��w
���Xx+7�|#�<�.�1q�E���*���y=2Th���0���oJ��u7QXW�.
	��FI��y���dE�A�?�j�u�X־ċ����Y��.ד�ﶄ�q�7���r%��QS}��
ɫ$gČ1y�И|��!
��z��wi���g���@��%���^��(��Έo��6�V��{;f�=Zq�� vw���ʥ]�**�u�W�3Xc��(�{0nފD��[�$}4��x�/����
���/I!4t`ף��U��/4K��˼���<hS���&�Yl����v+�I�}%����_�!�~�R�7r��n�b}/�ib�!Og�W�1��z�+8�Ȉ��lx�VH�UW��\Vc�F@K`1�Wx���� �S��Rp*ä�M�B���	T	��7~���T��܉zGL�ܩ�ѷ��(6��ogהo���'s�e�h�r)ߋ2+�6$B��|)'L��6�%��>�y���R:nxóA�ljԴ���%b'�/1}���;�-e��?b��T�A�`�U4�������v��a8s��Y��y��w#]�������of��|��������e-eh����2��IɖX�!��~�j0izÁh�ć.IH$(��W�elh�[M;�LQ�.�;�����W��!H��]#>'�=��h��eMpg|D+2b!/� )��MT�Ϝl��g=��a�I5}�1]X�_���4�<�:2�ٗ����GO�G��b�MjXX��+�`(]�L�mR�Q�8V����}���Eyy�d7kNF-!V�՛�N=���
�B��\;���<sCa�ԜUö��Z���x<�#�m� k����5���'a*a����G�T���E��vSQ0��	�HS���\��Q�$�D'h�Y��ā0��R��^�t�C�Iȸ���b,���ksLf+q ��Z��rW�z����1����D���N��mX�+�3Q��uf��jpZ:��Z��*(�%�W��t�Y��
�L�%����~��L����w�ti��M, �Uyhb�A��Hz��Z�~_%՟iCI�`YQ�ro"e�N��[^[�p����"
�fǥ�%*$ivM"��0�����u2=��X�2b�v���f������E�w�hV�<vKQ���s�m� �Z��ï��٘F {e�#������@��n� ����s�@��0 vϲ��r�)�>o�`v�B�i$aW�����d�t����	Ԫ�jͯT_�m��
f�␺x�N�F��:r�hq���I�ޛK�oDSyY��-"�T%�'�!�7���d�烜�<�i$��<8���#����F����qgD>R�]�����yp[��y��c��K�`T�������{�T�w��v��L8�;!��+�)w����͎ԃ{J����F	�a�ʌ�onXZ��Ŕ�dd8D[�(�).���qM�8�v&tԻ8 V�U@޽�#�:[Ｙ:�1�����/���m#ʎ��j>��ʟ�VT�Sg�B�ƱdwI�޴���G�w�i㘞n�%M�ǆ�0s?Y6���ue)�jٗ�8��s����~c�/�O�	]7�5MN����,�ز`$Hh�������6=��D���=�����ܓ�/C����|���[�c�>�h�Ҿ��>W����I��l�h�'��?'"���R�S$����56j;7f��SN�_�yh�����.�,�6���;����Xq
�ż.��8ʱb�~�S
ׁ�=�*��Kv���xh�m6K��q���#���U�^%J�����VJ�&�IW�:z��Tբ!���7�mb��S~�����(_�b��Rt��
��]�OͰ4{s�G>2���p�3��aV����U��c�w����>r�5��_ـ�����s.x����j�B���ϙ���q뎖��Q�#��2�K��!~�yH1�U�
��X/)�%�^BQ��s��HIT9IW�����	ζ-y����\N'M���2�:�N���{�<о -lb�xֽ�:Bw4�/��&`���K���g�y z�;�S���3��v~���^�x�����	fP��Ţ����-ٲ굽85k���V��	O�)��8��/Q��a����U�0A�?�E�p9�����y�j�|����?>�� ��a7�,��.S��3����:^��3���o�A��ؒ�l~�т����|n�3�b�����#4wL|kbi�܊7?:��|�e�k�~94"g�[i�[�X�/9��H�����U,����9�N&���[�/U5]��ԁGI&{e��a������2N�im���,,��\.(E4�aB������)�?D�d�˂��\��}7�(s��~�n���m�,��sL���[���"&�?�MP��q����.�����^z�`�zR�4��e���FJ]��[��"��.��94l5���>�A���3�b[[�[�AK�-_�L�N�����8��b[=��F`��U�pꑬ�1h�k�����L�,�)�z�T�<(�7�2�����%uon�Y����i�|���C�{�asC����;2)4�;�B�;m�G�nD���H����|�㨟�}�~�J=ˣ�Ұn������b*ng���I�ŀ�>�������3g7Q��u4�b0��K�gv�u%r�&�+��j-�v�f�$|���2;���]����OH��kޛ|G� �?���A��"�ʐ�IH��2i�7 ���X+`�JQ�_�t�Drc{Ş�*�}� ^���[�Ԯ��	�rߥ���u������+�E�;��	/s��й٦�����6l �Pw)���o�jG�b03�Q>ER=ff�jל����޴�$5r���Ά�+܏�sz���1Q���0�d���]�b����T#�[�w��/�G.�A<�"��c��Z�S!�� (�p���u��ζU�{	y�ʰ��l���LC�y���3X\�1�]�-�{'�Bo��^\Ȫ��ЕN�T�מ���t�0,��E���Ҽ����D�H�C�oͱjb���������)���p����^yi$�{˕�k�u�NU?��}�Y���*�G�7���_�̪��ge�r0M2v�H�U�
�����6]S�|a8�7�^.��5
R�l���}M�ҩ�͚~@�V�]���<�Pp�bu��>��1���H�\ޅ�MZ�Py��}��h����~	.C	e��Nt�׽�o:<\Αmvfb�ra���M�fj;��Z�c.2��pg����N�I��*~��<b�P���0?>�\[1?H��;�/����&��J���=���7�_L=o��^{뚪|��I��]��=�QG.39S-ǧ��eJG����|�t}�{/|Zw�";4WkpkT[t���ll����)x�C�����u���-�>e�Vѧ3<�j�B&x�ņ&}o�4�5�� �E��M�9�%/Q2�ȏڴ�� �mt����X���Y�>c��9$���	l/���V�\�NV���^r5Q8ODmaѲ�|����of1ג�N�����i<��F{Rc��ykS8�_�c�)=��`�����6����X6��%��C�bA0�y��IL�M��gS�%0�jX�W	�d�uk�T�y��Ͽ��~�"%E/b7[:$ٴ�,-��e���p�*p���N�,�P9�ژdK"Tl�7/=c�٪`�����3�����CJM	�WC�%e���n#��@���l&���vNZW~/?j���j����3ƭ4"I���
�劣;OE��#�����1�T��q���1MvB�������5NHK
�'4ˆ�a�����(wN�*l���z��K2;�,�q�����p3|����$UB�0�����k�=��VF��<�}�Z�z��1/�R��4���ƾf���l�YC����[���Z����%�9�Am�bه����Vp�(��ľ���a/���u!I���\s��U)��/���=����m���8�S��+E���~%����į�
���>��Qj�Rm#�U6�KY�����[�0{#�`a ���rk_��;O|[ć2(���#���"��lk����^˵h,���-�*7 �FW��T�5�P���N��L�ؚV�$(���0���6rW�_ڮ�����c?A�L�n�\G.�G$�,��:b����3A-��uo8��F��U@��(�P��v ��p�GyA�Д��r�p���k��X��@��e��߃��`wS�{�b�����운���d{V#Jκ(�-�͎'���/��zd��Q�8"����Y�OA�ƛ����l���Ft�W��0=�>�W�k�hO�)7m�^6Pw@߿rڤ$�K�a��O�SDFD�qO����n�sMK�)�6�6E]x��H�bM�gяNL�/S��1�J��t#�\H-Fa�i�y�ЗaW�5�sO��#��ʃ�>��u	�-W^;�фv�T���"�Z��$�> 7x/~�t����<�=e����PvW��g�8�Ƹ��e��v��)���W�����3n[����0O���)MW�|�$ҍ���o�N�)l��)����2�����Z����3�)�R&�T��3U�ƅ�%�������3�c-�R���ez��2�f|����Q���;�\bt}\Cf�c$w{��-rL(}P�^q������?��[���=����mg;�8$���(���W"�ui�p ���E�C�2�}�wSa	=o����.�����h�~:� w�ʰ���Su6�ery�GRE�WKj儯>���?�Of�T�{�ѽ�S5Z}�0zp����k�'�*���:"�(bt��r"7֔Nx	�1H�~5�gpnǓ����l���,I-�bLo� ڨ1N��
���NX�_5��Ҷj2Z�>�	�U��CI^8)|S��s~\���
b�<� '@�w-:��q- �f�.��*%�P;˽IE[۶PNl�i#B`II¦��+��*��p"�5��]�˕�U�TOV�rJ�,�z������u�0A|�j��N+�>(��+|ȝ��2�p	�/Z�>��-���������n���F`�}ބ��%�!dt���X3��Ϣo�w��\6RD��p�Oj��c37��<r��T�0���B-�:�jˁ8~)bD�����h>���C�G����P��rόf��P���9	`��[�K�d��<�ud���P>���_�%u�o�O���G��z�?��l��>9?}j5�����꿜g䗥u��A^��$�2r��o�]ac3|0���:�}�rU����8�Ni<�k��nz"�H��G����Ȟ�l������K� ��e�x���4@��|�
xZxH�}��dǍ��h�a�bj���PO�['g���#Ht�%�>q3
�������^"Mk7�8CǬ��|#e{��Ҝ�llN˓3`hq����g��M�9��?.P(TR���5ʣ�6���?��_��.<������pCE��o����&ߗ}��2V����U���^����&�v:�uCKm�8�����ۂ�u���s3�|>}�'���Aid�_��,sC� �D���X�q���B���96�k�/`��=���<q>��d+�VqZX������g)��FW�T�C�p�*�;��80Z4qz~���v<�&�y�s�H9�3�?�K�#XH�_&�9zrj����Z<�������e����d�z y��hǠ?� 臔��
^B�鹫3��{��r��W���&jG�8��\��ܛ�^��#�9a�>�]�9���~����֏�+���Ң��S�N�� M�����~��j��Z�r�0�ex=�vd�F�3J&��diA�E�N��hA� s;�@������k_1n��\���]w.��8�C	�[�',B�~�Ox<S�d���������/49]I�$�N����|ͬ���t� &�<=�.����v���`�["�/������CeG�h"!z���I�a�d����6UV�$�?�Ls���sj=`7s�6X��ݑ�ӯ��ΖV�����o���(��M�ɇ^k_�rd+>T�3t�,�����p.:  ��x�%u&hB�՛&2��M<O���<QAy���'�P��)g�<>ϫQ�򀤩ݔ�����d������;�=�F���oh���r��EY���ǣz&�� 71���-{��q�ޝ��;�VP�6�����n���Rs�ч�}��@Y��~��V3��)+}�'�0
�-=�&�Ǝ̀r�ǔ#}�;U7+�b��|����'R3��03郁oQ:U��pw)�����o��s�$�'~v��k�Oٟ[���r����$�
]�tȼ���j)��U�ؕ��~�i��F��|3����	�y���Yx-@�a����[e���_�P���+�����r �Gt ε�۸'�)��1�^aT4��fT���Y�����
�b���(0(ݧ{�nD��p7��ľ~�0��QN;_f��QC����F[�uL���F=�ZM|�
I+�M������o&�=BqN�1����`4��_�ζ�y$c*�+o�#���� �`7͘���,��o�>���κ�\ҟ�P+�2�L�)�uCV~'j��M�V����&-n6��@� ��6�xjޔiKπR����>H�(J��=scNe2L�1�s$�kY�`3�Kv�*�J����z�7�<�p˄���|y� ���Wz*Lw6<`��{ 	�1Q0#����}�]u��!˛\�F�l�k]�V��'/=�0��c>�+�*Z|�Ȧ!�3�߯�V9����ĭNi��u$�-��,��,
�W�+���}��x2�C�f�fR
/��� u��z<ȌK9>�c����3)�2�������0S���?����Ѵ�jC�ꠝm���u=�ޙ���j"5L����c8P���OO�����������k/�
�E�~TA�k:U�i5
Y��nL�V��[�����υhZ�n���!GV���xԭ��8%AG�[�;��-��$��~gAPG�^���%���J2�s�|�x�����e�-��|�e�xC�[��{���G*/��#�}��]xqj|H��7б�/t׹.yy<��<��߆��r��Q��a}�E��5�σ����Q��"z�L�$X��&�a��];΢����dZ���g
�t&5����WBy4�0g�-��M���;�+�+4ȅ�n����}�E�pھ�����7�k�M�C�;ΤӦ���0�"��{z�N&9�� ��p�,g�8ߪJꢀ_}��tu��W�l�ryU���"Lc�/0����m'�p+Ɔ�����/3MI��;>'����)O`T ���|M'HV�i�h`@%t��:���u�%?��"xs0/ *]����xrN��-U6� #o\4���j���/P���Y�;ש���;C�q��w�Jgdz>��=�;�%_?|2DE�T�>�Cz�Y.3���Ч�<�!�u�~�ʤ��P|��3��3��ͩ��N�=��U�H=�Ζ	�S�6�s��ze_e5�j��7���A���*y�[ԉ�(�!d�1�w�ѧ���ި��F2Ը�K'Ĭ������m(��Y�[uQ���+_����0����W�9�o6 ��"�p�����`��j#eZT�ɺpp�UZ6R�<^����vn���H,�㒒�&肅��D�&2\'��%b�R��~'��t�q����?���[ �얲��Iα}�d]���姠�7V�����cM�	?��|���Q̫�)�Ns��J �lU��,����ZI�̖��M5A��>�� �dj�d�LH^x�� �m�?�};��8St����6'9�>��Pk�m��^]l���ޡ�7��d��nD2}�]�`C>�̑�ݜ���_�DF����O�\Q,#CO�����'�0��kK�ܨ9<�?���0󨛣ۉ�8U"ߡ����ld���G�W�U����KN:��̵[��I�#�$��P��q�9)�Z�����6��9�.1�y�Fx���ȉ����q��L�k��7ậ��y�C�9�33-��^m�!Zi+W�J�CU��py�(���#+g ��6ҵI��U�S�/z�\`�(2M�������Np�GX}T����tw�"�P��B�]|�i��g��Nt9�jm�TWd�HvY�}������T1�q֢�M���G���	�DY��S�蛿jl�go���xƩgQ���(d5�����=)���s/�>n&A��hwn�̆�)e|Z�F�#��`�F�ܐʘ�De���]�)q�<фE_)�������LJ�f��B���=DėIC4Q�������������<U!;�p�X���_ p����>ٔ�d%ΐqfAгvW$[�_$�����F�3d�)]�Sk����0���
_d�r�s/�aDp��I��p�IU)x��>���U:v���kNRB�B�Bmh!���j��H�*!?���V��N��u��*R��ˈ�R�iF�qZ4�D�j������)k�էK4+QG�m�3�ͥ���������x�$/��Y�8��=3���J���;W,7��B��=�x2g���
{�5L\�*^�ud��hD��?��.Q=�o^[�^*�wA��.Rچ'�c���wN�CWt�R���S�e�K�
�˒������.�b2�|��|�E�?�?��d�GlùDd�ËĪ��=��+L�İ_B)�ʊG�47:�lVk��{�=�Zx9����+5��.y&��+^�!���a"Ǧ�|��Y� ���d��7���c�)t������9-���=����j���)B��y�o5E�B'����EӘ��R:Y<�7^�W����j���3��C�s`��Dd��;(�,Ӧy��Ǝ�U�w�Άh�ֻtO�j�e�0�rP=T���݈��ko����Q;� '��Cr무i�2�͚��] ��6s`R-�-�1)�����#�E�� �A+���<�
"ڪie}�A����µ��:f����s�D�uj�/j�LC�U;���أa��A��+����:=�%�K��x�*翢����?m�8�k�YgΉ���[�4��A��)1�**���;~H��m�C?�������"d�,�7��d���'߫t��N]�������;i�\�R?��U�7?Y'0KI����:B��c�k��ـX�{���k���b�C�#����ٲ�i�Apo��.��YV��ӀF�� ��3�b�l��z��?�1	cB ���"���<�̰��+kgٿ[���
�
ZA�35�LZ�\�#c�	�k�,�
/hY8�k�R����7i�8H�M�+�������<mg�\5s�g��Ts012��.�pb��hAR�i��ث(Ym)��ܖ����,?wB���^�V��޸=�>?8䥘���`lHg� c'l�G����������1�|=�Q�a���>wr
���9�����}MZvB5��-b��D����Ɨ}"ԗ�[xI&sV+pk���Q�M@�#�1���1��e�kKT�x�f�Ή�a��k�>u3��!�v%���Egh����k
�7�[r����.��m���9� ����tsy��_�|�W&�@�8��|���rj	�'���߻A\}���x��r��q���-���2+s��}�l��Í�!Ll�ecA�+��X�1�OO�r��YD�lS���V���Ae����
0{���G�(��f sp�������-0�OH^��_g�:v���f�:�3��ֻ�V,f��wp����1H�`�ݜ�#����F�Z���b��ĺd{t���sN؜s�o�+t����,�+��(.A���� {0�4A'S��!F2�o�7n��� ��<���=CJ���r�v�= �>g����P�JYsٸ�1P@a7������I^P��Ӟ�� �T��jHf�{hw�<�Ԏ�� PKRu��G�{�V氊J�Uzn���[(M@�\�U9����L�8�A�.��I��|vU�F:?��;J� #a�O2���_a�rR;i0�l����[A��(��?��^g�)��n�&y�g��j�x2\X(t�x������P���&�)�}~s�}��0Py>=$Lr��@�����>nE��f�bK��!���h���z�����e�^!"��g>ӳn��O�V>��7K�=���x�Ä�Z����a׍n�q6�z�/�&�V��MG��G�Tb`Bͭ��w1&�:�Ϥ�-֫�͠�KP��?��t�v�7�%��t]>����1%+)ьN�ˡ��4�����	����	�o˧����s�!E��bպ�qR�L��e@,�M�7�g������0O(��_���~�V���\[���jq�\�c%y��ũ��!���Ja7��SK�̍E��!���{�<���EyH��EhW�_3�b��F��銧ho6e��6 0�qC�x�ˊ���/1U�ס.�m�-�fh��3=��P�N,���2���%�!��}.�]�WK/�t�i�P���i^u&�mosx��S�D���r�����'O:�J���x��5�"�r�c����� �M���9Я��*�Ƙ��x�O�C�Y��@�\Sc5u'o2���B��n�y[f�y�K�$���
��2,$Z+��h38l�G�ʜ����`�}�~�osH;����o�iVI�OW)F���Y}�[W")���GMQXN�O�ޡ��Yh�0+��������&��,#Bv��Q��V�~w�P-��{J�ʛ"�]���|m}�l[2�T�3�W%:!��ꗓ�r*D�y�:-G��J��ۚ���}}i�;pKx�����⼭��{APPU6�7#�S�ǒ�Q�x�L8�5���~�7;�ʌ!м�@37�-!�� �/K�+��4�O�,��*��u��+��-����[17�xPp�%��8���2y��O���#p4�<�x:�h+��lǠ�.+o�d�,�v��0�j^��9�bN��v�G�[������Zё���HF-!}����א��D�|�o���F��XF�5���nH�Δ��MwU)L��lS]�U#�	|�-�<nӏ*�Po��̎�-�OtE^�"�ܱ��IIyNz�r�����X.C�4���g�Y΍����k=�Bn��l��04/�.��g����~[�k�2�̾�e��_*�:��r���'��jNQU,��0LD@B��_G-�01����ϊU3|����y2|��$�U���);����M7�/�_O���N��şe|���;R0|w������,��5vs�VD�D��T�6�\u����ҀB�L���E�����mZE��A2{�l�)2~3��Pt�1|�hwP��Ϊ?@V�IJ�\��l<3i
��E;AV�,�d�NB���^�����LX�fH)]�t4b�|
���0PYb	CZ���̲����.2@C��v�ǽ]L�l��E�h��^�`�.J�W�I��쪩bmօ	?���I�.�q��i�D��fɵm��Z�Ul4c�n�tx�\r���(����q�,.0r�Tm��W��r���>g�JPG�j���J?E�i�B�d˴�zA`
Y]�$fb�ǿ����+M����3Q�T��'tP�#�uP���K����!	�O�⤁�%]�a�f5���������^���SsUL�S���*����ц���PS��7��11蒔��L�����[c��+���ٱ��H�w g5LD��@ȏ���Q}��L����Ȫ-��ml�pF�sk��F0�h�\�0d����<�E�;^a��}]	M!��"z�/4%�6\���$a�q�BrWѪ���Z�uF�ce8((bi���=�+!��T�����jGF�u�6�g��Sl9n+�:P�v��fQ���u���80��Q�Л�ƈ���GYm��K�V��b�
�is>ɛ/��A�U��������2��υ�PUD񰏱��r5��c�+� 0oNi]$�%ixd�l���4_�㝫)��؝���`G�|L�%����Z�r�lnqw1����F���PIe��ׇ�?W2���^�7�`^;�������[�c>L^�*'�j71��Vtl�ug.�ȦJ	?:�w�C����4F�	�-S�̩@Lw'5l��CYԡsOV��7?(Ne���_
OA;���#�,�9�`�egq�r�C�4FB�����&�p�%'�,ۣ�����P��D`�����k�l��*L vӒL�(I,ra�q��;�l���#���7��9��P�G�%�@kޔ�g$u�[��)3̐ +E��B2�����$cRa�w�M't��e�C�����0�~�\�������[��C� (߬�Ÿ�������]3�",j���vҪ���������}qѫ�����~ku{�h����y�HI�휪dW�-Dּ�
̄ޔ5�(�`41��l���]p@�P�1؈�/�CJs�]E���>q~ �0���9��~�-31�F�f4���hh%���,*��}��:!�KNm<�%�h�����ddϰ8_��͜�^3�H �����`�>�>l��C�8�t�h��7��ʁ�l��p�S(F*�:���~�f��|�gs��B9�D�`���8O �W��XY��L>�r��v�gl�0E
<�]�S	x)�v3�I�uЇ,)�lJ�T7��̓�0.5M;��̹N;�0AuuGMv���}26œw�K�-h2`�3�[�V�E'Ѽ��@��-Ѥ7e�%t]�3�XN���4����Ȝ#�	e����]w���Mn��w����ӳ�@'�r�zt����ږז,t}]�E�)Nh�Q�`��4���J����V�`�y�)�~d �T�cH���6�'Z�4���SO�n�*��Đ���8?�S�@�GN�+��}�C�(��I_��Dҏ��l
�K"(��Iq�uDTl�N�����N�}0Η������U٨ph�d�cZq������+?�1��{���L
~�n2)JK6��9�'�5�u�=��j������+LY�!*!Q^s�ʥ7#�|�����K¶�@��n��+�g_9滴���"�O�v�	+m�zϥ�f��f�z�"^c�����<&�x(t�C�'7���2[& ��J��'}\�"a��v�g~9��1m�|z��m��üJ<X����x��y��]�Z�)�6`*'_q��pe+ưW�>�Ԧ��FE���S�J�3����Sj�x���A��?��ՉnI~[]�yS�8#~�;%C�/t�ЉF��x��W�ǿ�X# ,ssA�ٓ<o��j�l����o���gIo�X����&DtD���e�#AP�ʀ�d<�Li))Z쯴w��AqJ����^����9�@Ӛ���+o3��;����&\��/���B<������&��0�<��ܮ.r�C�&b��1�8��}<�0��G��"�� �"�(�i����C�ە���oA$,g��Аk)a �d�P���7=5�!�/���q������r:S�����?��`�e�Iorwd,���b��1-���]��md���uٶ�JhQ�nG�A�����~Z��'��k&Y�cY���O���*�6��/��oU��z�g?�c_W5�lde<�yU(T5�<5�9���iu��'��3�PгN}��zv-�e���iH��
= ж�:G.@���Ofb�����2��ǽ�(�N�7�Τd&h��0Zh�y�n�E��e�h@����O5���>�U�Y��� ���Ȋ��#���m9��C,=�]6pit!T��{��R�~�L����}��ĶȀ� 
#x`���7w����Fq�Pdʷ��V�s�M�&(Ύ�F-UF��"��8:��_t���F��e�.A���խn])�r�Ff�kWh�z�;���'_(��3i��|&|.��M�*�_�9U<o׶ ��n��Yia�c���`�9�����bv����;~w��sƿ�IZBł%"[���J���йF�x]-o�J�J��D]��d�G���߹�A��gj��ӆ���	��s�Jiq$�M��N���𕍶-�0/��Ѷ+� +��������f.�L�z)6*߉QL4��C� !�! �
�k�Cً�ʱ�&��8+��ƫ|cj��d�6c/�4�ʬ���9��OpK:�y�������cz^�
٦:V.)�������<��'��f�8[߬��d���� �w<���hPӕB�o�c��#��3�/]/�55`��h�]XѷS2���U��ᨄfaP�x��=�I����@^=�`y����z��]��<�8?��,�ֿA.�"�U���d�/�j���+��?���Cf��m��ኋ����-�{�!:Vݺ'Z� Y�<��6�`�r���_7��U����&�����m[�HiD�2EԱ�Yy�+S�
��~��X�-=���i3�j���ռ�>�B��	8�BX�����k�9���P�S�� v۴9�sU���_����nZz�:��V{��?R��$�Qn^�����z�H���R4�N�6@`6���:�bVVA�1?/ϰp�*f ���km ;+x�Z��\K�>!����h3J8WC�˔>*�ne�=�c��w��\3��V���Xi���xq/�R/��VP����G�9�:��*62�X�\9�ͯ�� �[��MY����5�*A��D��a��y��H�!?o�#ִ���d������>�1~1�!{�X��hx!�81Į�����Mǵ�+�O����}����/n����7(���5������Jf��f��g@��>�f����թae	�?[R�;�C�]e�]D��]��=TJ�U�h�!�M��Qﶨ(�k.t�C�[��C8(��L2)��D�͍��xR�}`���c�!�C��T&r�tU�,noJ��m�R����'F&��v����7;�Ww�ɛ�ئ)�F�¦���fݷ&��n�U�`G�����Lb�ϐķ�?V��Z����y��k� gb���,������u��m0�׫����M,�!`�	E�,&��^B�~�?v >�������[g4J�Hz_3�������QС �SI��/J+���Ͽ=m݁)QEٓ��*�'���%V4�|����؉��p�x��Ш�-�����z�:���AF�D��0�̃�A��2�ݮ���T��d��� ��_m�Xl�Ш��U��w���pI`��w	���a��݆`�S�A<��@�#&0��i�Ra6%�+���C�g!�{��k����B<I^�Q���p%i�;�"�~I�6K��8���k�D1:9C<ݗV��e��tG�"�`��E��kXS� ��&�z&�H����
��c����ЩЎI
`ߺ{���^�]��~88{�g�Wſ������F��]�ý_я�j�"z;�dy0�`�4��0�W�j�;� ��:zم�Zh�A���p�?�{����Z
���or0T[����ǥʘ��i��c�Ԓ8K��iL;RZZ��*��K<~�N�AA�mM��
e�c����FkVA҂��l�t�������X�*�	��Tr�laq�v���G�iNAt���ܽ�ʷL+����#@W�L|���_x1E��q��4����]Z|�Dki.Y.w��m��>c��X���Hq*$+xK/�y�q��/�����"@jo8=�N{ɲ$?j�RY�ꂚ��)E�@��애���Ů,�c�q�T@;IO��c�D�#�-�-	>���+��] ���>D!};��:)X�����M�-�#\j���3=�6��GW<�~���ӝ�wÅY(?����{�q�ئ�:�e>����E8���3����=Z�{#�n�jk�n�9�Ǵ6&�+i5j�[؂	ϤI��F���#�����$��O�V���W�:GJU�>��0|?K��w[�Sń������*��4/N��"׹��|Wp�f�(��FU�~��;�5b�6��\]�Ao�<Xj{�Q�毛7��ՌCO�:�1i��Y���z8@�����D-��5T#��݃`����ލ ���Lm�%�%Ip0�x�sٚF�����Ik�ԟuּ��LH���v@d���J"��s	'=���@�-�,ǆ��B�k�%�AR$�[�Pd&`0=�i���*��8}� 6��������r ��c�L�g�/`r�Y�V����x#�q��ѷ�ժ^��
{��H?z =]�nP���>-�_A�9��\B�*�%�R�� �	������ln؊�r �%agW���y��Jȿ���6Yy{l�/����z�(�e(���V� q�*�����/i\��K*�,�\�V�����IP�Pzyǟ�׎\!�*+a��c4Hm�#-�e{
4j7�.g��<���y��~��o����3�b�8�e��ޔ@f�Dl@=�o��u#��_�7O��� ��N�`��̼��^��@����bN��''-���7I�ɘ�WU<`����S�2�w�=WGR1{��U�.�0B\��`�N+��FZ.z�M`<Щa2@2�U��>8��� 23%8>D�����l�����[��HS����ͳ{��2�(�zpb����� �S�����#rH�z@��k=YNefiF��(���������]V7��"	p��5�o:�M�ʃ'/m>�^��y}�/���sIK�lB��	<C3�<�,�,���kD|Ns��i�]\+_9�҄�V��t���jF�1�*�׺�p��m����xKI-��̷4��Ux�\;���l��z�����+��1�%E
GQ{EF����?"m�q���,���R;@poЭ��3�� '�}{Z���\]��S�[A��α�?�=fˎ3�|qq����ά	��.���#-�����Ψ�|w��oe�-!� R�2��Hk���/"2�#��a-Utu��ɱ��o��5�A|�� J��Ll�[�7����m�ץ@N���L`���]7��t��BDo��΋���!	.K�"�,륷)<���	w�����+��sTP���tc �S��lJ����ڙN፻|�c8>*��L�$���IGi�8��&(C~7���JJ�+A2��0?��C�$<�9Su����2� ���xL�t����?!��b�b�{s$?$��]�jx؞���Nvzk�	��◙�DP	���!��_�{�����~|�Kڃ��MA�0���uJ�"��ϮoD���"�V�7}%�X�d_.���`K�`,�D*I�x����� Z\�檃�g�ɩ#����-'X9ʤ����du�s�3I��(��!���)�q�+�������f,��U��	Кyf⏶�mot��SǦ>P�q�^M��D�� �|����H]�g0C�t��?C���|)_$ju�-�1]{0<�~HM�z�FW��Z<�)d#E^5b���!}�1��}H�/��}������"�j�1u��U�R\w)�k��-v�D��<�SD�����
�zmg�2�~Nl���3&�B������e.D���8�v�ZT M����d��%�����n�*�����{���/�_���$h��5Y���?g�,�P����F�U�0�Gb��k�}W[��I��K�R��H��]y��yj���{�RL���QAPi@A��Ő��U${!�*�pu�6ZY �e8�A䒹� ���Քu�A��h����83�x��!F��_,����ȕ�[X�_�;6O������jbt��w�FG��jӨz1]\�Ҷi�C�%����P�Ӕ�{Q]}WG��j��/���	���83z�ғ���_�d����bd�hu-${hԼ�r\H�U�]���>fQ�n��T��ƃsdoC��.@ſ�t��ݙ��3��b	��ך%�g��k ���Ss�1:Dx2�V����L�K���q9��)_����ND"n�wu ��c߁�>�DC����['�����[a3.b�Pe�X�~������?sK�1�OPˊo9�";���s7�`^��jPP�nܵ�g�
�[ˣ�eSc$p���v�1>ð6Dò�h�9O�@Lj����q��H ��������`ف��_������)v����=f����F�=���JL���Ѥ�S���V��s�ss:MG[�k���s�&D����?�UL���P��k;��-)�I��ӸU�n�e�-'�"rF��9��Xϩ�I�S�4`j>�b���<���a��^ l��q�ϳ��Úat}�M�i�Ȩ�����맦��O�����)�W:�8��@�yRx�0FtO�y��4��>�x�������kSݰR��+#�DrS>����sT�[��F"g)L�x��f���MĠ� �$j,N�i�6�*tl}�]�a5������b�_�%�.`4|"+��}U���l��fKҕ�G<�M36f�������!�����3`��ث4�z1�l-�V��$L#���k	�v�����t�/9��c�}��͏;x��^u�M�Et���Ϳ�p���H���W�������:^n��phO��t�Z��A)u�ti-��K���e��TX� D����3�u�h���o�bYy	v#����� ��S����&A60(�ϳ������/��0�r� ��yÁ,�l�,ψ��hh>q@?!�-�E��
������J�<���k$t� p�>%����pʱ�r%5b8Pr�b,.��S��2��F���xM@l�@OSP�����`o�.�����S�S�������r���>�#C�
�2�Lzx��� T�u*�7r5TS�I��X�����g�kz�a�w	=�# $>կ�f�382̟�����κ��?�.���U�����J�g�8��hT�H�����Q%��1Iӕ\��U���~c�`5U�Q�T����O�	�W�t�?2���4y?)�u%I;ps3XW�_��A���6���֓��S�D��}�.k���uIЪԡ����g���¹��YG����2�Z�_�8s�=�t'+�~��+<��7Q�/���Cû�/�'�x�<m�Ǒ{�MugU�)��랬v�&�R*����~�����G�t���g$p6rh9F�xK��F�l�ꦿ,(����!�������ǈ�m���Jt�� ��-����:MvF$���v(w�S&",��&:�ɨ�]����;(�h�:CG���@]�"�u�V���\����F�%F濲�>%���EЗDB��ۥ�f�*�R�_��p�h��ݲa�v�U��:.��n�39�g�+�^��mO?�nh0�"��tݩ�9�PR��^mG1Hu��H������y媭U�>w�I��X�0f��V���DGcP8��ӦD5)���g�)ZD�^)�cI�/���O)С*�u2m*�bO�:�c�`�r�3V*�9L�wh��V�C-�Rl.�`�D���=�W�FO�����BnJ���,l%u���E���2[ь����&�e��:�Y���
V>��$hU6E��Ú,c�0�(k e4�7�r�%�NU'�X�M�T�25c�����"��HA8C��\ao����퉋��X�y��~?�T�4��0Z��0,h��˴#h�A��	VHjЖ��)��ңWJ�Z�Vd��:nK�U�q�#�&�=0|���79�[+�C��WN�E�}���p��6��sS�S�U'=��b�ʻ�v�9q޵���r]q�"P�� y�}~77(�F���)�ʟ��4IOo�J�|^l�,G�ک�K���phSW�&����A��Uh�S�&���5w]��w�m���t����S�C�|���� ��}��3��2U�i0��J΢0��c��Ә�ǚƄ/s��H\mnq6�0���E`2�ONl�g��{��kz����Cq��S-���Y��4�B��=�4�?�(PɁ����.u�[��)���C��5���8|[�x�6Q�W����D݊�
�����dy��:(I�#��ܖ��>E�ְ���ړL�r�%�F�2�
r*�߁�`Ǡ^͗
�K��E�G�b��:ԣ�ak���Rl���F�{HսC��=j�����Q���/Ze����ޯ�[�*n����Ne�Ǹw��E_w��'�6�+x�49�$��<�˽;�A��G6���ʏ��O �P�����i���b�I]9��$m��lc���Hs;Q9���8�����7?͠c\±��xd��
y�����8� 6����Ӫ S9���٘�ieY���g#�*c����.M���]JS}�(�����Q4���*�h�%Bڔ�f�NҠ{{?�(�#)՟����6�m�o\�c�� �A�i�7�3{l�XY
ng���R��C���U4&�8uF��.CG����ֱ���MkB�F��_���y'��MR��4��(�Wŵ�����k:�>�:~~��[|WYv�ݺV���� ~�c�V'7�@~�/���W�$(qm����h�D��G��MÙ�A��A�O�+S��`��[�}yyy`�����Ň�Nb4�vc,d��+�] )�9�W�ϑ�^�b< �w����o�
-���4�=�cuR��h �}�i����o�voGX��a2�([i��)x����?�B�u�`��Ҵx.݌�Ċp�����%�6C�������mlo�Z�%Q3�2&�h��x/B�"Tw�0����x�d�
r�v	���Z"Y�CZP%ij{4|N�	�M��B��Z���ׯ�x�]�9a��]��eabS(B���4lWZ���Oh�9�۸Wٶ˶����N{N�>��o>�]���_�p����ٓVz�c��p������w�h�D�:�fi>���0���VG��ܒ��1�{,Oj ��6��ZlM^������̰�?�ۺ@���T鹝!���-�������詫6�n@�ZA���?��@���;p/�}�y]�Ʒ���d_z���0 �a�h&m��?�q`�X����q����>�� �Pax�*cL�`\�i>��V	�L�,�9%�2m
Y-�����5r��I$.Pr�g$J����MЏ-}=M4��+n�{n1WW0�~�O�P��GL6���㺇��@��"��� c$��n�4Go0�r精x��2���M6��(GA����Mas eb@HPQ K�'�XC0ZP�-����BiP*�����	��x"����.c�=�'�Qk�����:���s�C
��52�����c�����Ў!��%1�]���.�CUI|�׿5���Y���	��I�� ��Q\��Sov�V$X:H��.�PR�}�$��$2�H��J�D8l:�؛'��]��r�O˲9Pj�/*9��@>,%)Kk]:�o<�W�5��	w���ңC������}�i���A�&M]]��#�:ј�H�-��2 ���)WP�3d���ʶxz�7��s�|�:H��nz����8�t�xZi�/�����qf��}�^��j��f�%���d&��F��%��o<ݒ��UQ �ڵ��@��W/G����q|q+��ǵ�h8-Z�U�}�j���ɷ��+$rӔ��ߖ���s+5�ao������D�8FL�3��mc��;g6���.����~?���E�$ZY�>�<ȷe~��-�.>'�B+w�6���o5�J&�S��is�ƘC��Ʊi���ʎ_a=~nީ�?t���D��vu�0*��1Gm������MXt��������j�fp�P��Ų�#ޫ�z���ѯnG�7W=c�c!g� �-���r����1��'�&�B�c�K9�>���������{�RHҁ���=(�C����18n�:)
w�޲R����2��l��,�ǻT4t�B-��j��J��(1�APk���u�V��F�r*�)����8Fa@o����XQ�|#������1������c-(���9ˍ�mm�
����_���P=;����g�O7��I	x�<gL�7��#�v�#}���.k���j6N���6����>�p{�v�r|�1�A�a,;��_'*��h o�-�)lg ˰�&���oa��!�P������!9�XV	K��R?�٠B�z�_��>�������������6�(��v|e K̊�*�5j���:���x2˙,�U��W�T�F_��Og�T�zM�Z���(�����3�����H�'XB��c㣜���M���&IM{�DY����]y�w�г��4��R�Uy0���?�d�Q:�'%9�k{�@��FtK�랟�{�����>�z@}&�;ݷ�%_��txv}5��14Z��秅a3�pW��$�'��{�tL�H��Z���V1�Y�6�*BM�Z�� ۷������8�wS�
�:�(x�z�@!I�rl���܇mEӹk��� ��b���:���B}#����DG���ei�'��o4oN��Vw��*��48og9����q�7����|��߅�%K�nOBo�2kt�y��X�<��M*V��a2������p��ZQ�Hd�w$8wN��[����m�v��Su�D�Cۨ&�U�	ۜg�#�c-?O�"V���i�eG9!t
�������� Њs%�0.�V[�dM��W��P���o��^�w�mɟ�h.���9��?;~mђ�Gkn��3�ZFAX��6���F�\t�:Wr>a��i�9��)�т6ᛂ��­H�͍�c�"LA�߼��ϳy�"5�Ó���W�
�
`��2���{U;��<'���8K���%��D�A!9�M��v���S�ͭ�=����*�;
��<��F"B��s�����~�k�JP�o��kV��4kՊB%�fw<P�o�HL����;&T�9���j����T���'�y��x�X6᪤DY��)��{����b�6�`lޏ�ý8����]�\m����l��H�#�����Ѽ`3f����@���^�A]~{�����*|��&�TY(��NMoU��P���/�!u�%"@�rݳ�u��[q���I�č��xS�PJ|ѧ��1�i�I}�U�nqڕ ���ݣ!��S����X݋���]���uӪ(e/����yL�y�ߠ�ML����$�]�c���d@�SH��/�Y��}�5������k��ɤ�l�7�0<��~ꁩ��;A� V_�/}��cO�W|������&Mf�Ǹk�J>S��<X���-)V�y$K�_�CN�H��P��*&\߈ cSn��������KY'_��V�hq�J��Fo]���~E�H?�dr^�w���E�e�.����mS9'��R␉�e�&�&���`)�ܗ���ep�������b�C�u�?��s�L!�iC���~�C��)����\8�n)oM�x��JE�'�y0ϻȥn]H�3�&=����qR����q��c
P�K�C���\����ᶯ���0MR�;�Z��,N�X�\��Cs���$�
�׽�βa_IjO�!+}�\_5f�v�:��y��؀ȁ~T� ��i�����vrG�S�}Y��~G�kҽ���ԧk�)p/�,I���5��E�"�M5�95��%hF�[
�����������&�AǓR���۩l�����pn"�����n��M9Zȧ�k�Q�� .����+��NDz�3�7�|S�Q�m��	E�F�Z$Y�R(�U.�JFo*#@�[����0����d>�׿�z����@�<�d�qX�,Ue�����U��'��Y�����U�)����n�S�4we�BWC6[���=�U"�#�����+p�ɥ��O�6Ӹ�Ѷ�3D䵢�J���nĲ�J�Aj�{�N����/~��g(q��1�q0�G�x������&��s��2��v�dL���u�8���~Z��bK���]�J6�Yi��*E� �Qi�H���^�f'	f��
f�����7��o��[g+���[܊������^շ�g���V:��4���f<�U67d��I�Y���y��]=�����<��Qr��?�	?]�*ل��ޕ��~�{�C�R,��n,-~:�A]E���c��ANʓ�H�V��<�Q�vlY*��!4А�Hi$�B�s�鈜��ô�{~��`نo�_R�L{�ӌ�!�l�# �p\��{x�����\L�eŀ8���{&o�8��|*�v�2���k�N>ՠ����!�ee->	�������-�Ur��S≹3nc�W�6�XNM���=�#'+R¼��r{G阗%���!D���dѦ�^�fY��&;wx�4}�6&���o��*�cL~�֌�-�j��z�%|��]�嘴K	Z���D�_|�W�ڷ��z�_L��'��E%�C��w̶k7�wS|��4wp�I���Z7�׻jq����6���g�	�b��� �9��*�g$~��z�AUJ��k
w��|���F%�;;�{�Ɂ]�p��d����L#�184'�b=�$%�<�O� 7�ܟ��-���߳=����挋_����ZД��n5s�[U���>!�^W������w}	�ȩG�[�#���Z�Ё�5y�$��wr��lmb��z���\�n��7��]���&O���3�GV�MxZ%��X�\La+�s�LX��< ����hi�
5�X�20v�E�ڴ]����N��x��C���������k��!�����������#�l�����١�/$)m7/ �Ъ+DW?������	2��ǋ�1i�X^��7�]�^Y4�8 �6�����)8Ԯ�wҨ��7c���^�	��Q��ى�Y��"��dA<3p`F��%�%s'�,��&L�:�ac6SFWf&\b�#Z,�ȥ�/�KY�E�h�?TSS�U�yUU=߾�hW}�σ��"�e1���S�&�χG_���1=:�>c<���l�a*�f�8-]�ڸ��s��T�^�4?�4�vw��Z�h��¢���N�k��3U+�u�7 ��a�~�ur\�:㐩MR����8�X���VA��@�Ƭބ��j|w���] ���ĵvyC�ח����~�zI�#P`\Em_�L��9��+��8R�����O�x7y,F���H,菉[�����$�}��8l�cY�ͷ���l�A=lB��a�o8U��u[i�O�ئ�+�i/����4W�tħMe.�����]w`�����U��>ўJ>��B���2�$� �1��r��d|������B</�ӊy�ϰ��	q�o%i��	l�J�3��1,�T�P�QY�/��+���"�(\	k�O�Ҽ��mw<q��u�_�����4�/�2��iՉ�R���@���ݘ��}�s�N�+<������8Nz��0Q�x&̵��&�:Y=���C�p�4ZS��ꡞa�m7����2�z���7,~�}h�����{�C�sf��+���z*�*+��q�k7}b�C��r��B��;����T�ahE*� ��RL��֤,�v8�ȹ��l� �=v�Z�o���IZ8a�l�F�B=�� �i�<l��� �:W�jl�-������}�~ؖ��ahI�C���4E�����E¤b���v�)^/��m���M�D���R�v���0_��0�:�2�:�7\�]ó�L��-��_g ΩB���%k7�nI��}��+7����˾}�H��S8�k���0���p�X��} ��K�6��l(����#�y�'[��*P��P�̷v11|�Ծf���w�V��� �@? �*-Gi�}\�Ub3V�l�����0$��<Yt�E]<� �e0��ioEz�	�ar,_R�u	����ua��^&y#~�z��{�3�^%*Lס>�O�]EU�J�l�Vj{�N��OF��n�!7���f�چ��6�]�ʦ�q��U���4�X�(�G�
�s��st8�������ܫ�|QE���X�K�1g�6Nި&��=�u%A.wΦ#���n�~1��m�U��欶��%�=	p�q��L�Ώz���ƣKv���7p���ޞ�
���~�ޅ��G�q�n�D+�y�B5�4�k=�&��$��:������o�~A�H&	��?�u	}C}�bք�t?dw$�1�IJ��8�;fI��>�.��?o�A�`2@Me��L���)UMB	�ު�g����~�A	��3�4W� ^h��ܹ������T��a��y�r���������',^���'B�T@��y7���a[������[�7���W��'3W�7u1h`'FX�(]@Fz�d���QC��_���1]�oĚ<4G3��W��U��������@������3K��To"'��?�{^��m��\��<o5��K�t����Я�#`ݼ5��1��9S#x�Uz.iz  [��n�]�2�sH1+���8y�D9����&oY���ۥ������Z�'�Lo�ܞ�f���hBO�2�J5/@l�&���r�㘮J�gE�2\Ώ�$��ۻ�_�q`��3��_��	
�1�X��*��gW!��~�����[g	�t(�����d�j�^f[����i���M�<��X�P�8e
�H�E�۲�|�#�)��˪����Wa*4��
�V������{�R7j�~XG:�a�e���d�N�,��Ti<�u>�K@�������/G4�@�|:ƶ�q���8w��Z�Ck�괎�^��q�87�͠o2ԛ��(Q�������A�.���Ky�+��vM7��P^z�Bl�Ԁ1�&,>Xs�:�>��8'��g(8��( ��)@�i�_6~r8#�u�$�nTy�}1`�X�_���b�!�:l�WM�O�k���3y(XҊ��j���]dp&Q�,¦��s�w/� �
_	���NҴ��L��	��bE�h�Z��\(˙�5U���j�vcET�p�aү7�+4Y ��((�l��+,ѓw(2��P&�0t.��T�o�o�!�9�u�Q��&p����^	}g����ɮV��Kg<peH�����M3м'�ݯ��GG�~���O���ٙ�N#��6�!�C����V�%ݣ�r!j�-�N��,�wM#�ս,�4�Q��WFB�.����߾������am�|�
�M7"��A�,VW��95�u��U�K%uJ��D��Bi��_4-Kj���/�`�2���QRY���9!5a�Ɗ�� *ߑ9Y �1v�L0�r�*��;׬�	���#I��S)�%�}�{�ݦ���t]2��ވg���G_�1� �Y�[�d��I7)۰�B��!�F+��(S`y��H�F�
˟�Kn�:O1����N>��n���u�2=M�KUP+�����aM�ʒCm�����e���M�	�(,W�j=��85�����i)pxNMi�4}1/�DyԌ�d�	S_R�R�D����{y�l��Tz��7��d�7Dg�͸���5/ʟ��c'.�?������|l̪��\�������@N=^�{{�xA(����Wm���DךO#��xI\�i�Vr_F�E_Y� �^�;r�L��*l� s�3x��m�QyQj+�o�����{�4vY]`�K�6=RVe�����Q|�J�⺊`�+h(�7G����/,��Y��]����c�������nTk�Df,��|�e���We�4ң9a1c6J����ج��
�͒�t��q|��ڽ�]��v��im�s�ϑg�����AbIׂ��w��985�]5�rs������=�"r۶�Vސd�=��Q/���N��&rH79�	�y�H;�Y���~��&��+���/MW��H��I�Ӝ����a��US�M$Ԩ k��OD���[��&�D����#��G�c����C�iuØ���$)/u�0 ��s'�y"��h�����f�̫��\�u��Xn��k�pz]p2��Ѓ͗� :�:�; ��6���m�*a<�M|��m��Fhja;C�\u�%�uw��6�c����Pv% #F+ǻ� �Y����h�ȑ���gE�����I���y����Pl6DJA ]�q�)���������m	�m��1�3�ŀ��I�����S�� �)����@����6 B��qv�&N�}�A��i~=�c�BZ��$�b|�A!Dշ7y�p����']�r [����W��b\v��(`5FGkX3��ɱ��II$W)�Y��gm�;��2�@��(�lt�?��t��ʘ}ã̡v���!�?)�����R�{�4�Bڍw��	lE����O�X����ٮ�d�흈rS��-�>�{���R�0Q!�����$���+"�	s{֞J릙���lv�S�Ja&�`c�SdL�P@T�xT�������=�#���E�-��i��[��2-R���&��c_I����9��s��&۫�.Y�*)ץvaj�59�t*���6��ަ��Pʻv�9�s7�YT���KZ�$Lg�PsE/�D�|nVv�u\pˡ��,�GP�Csd����w�n�b�w(�[�
���[@��3e5���ۓ\b�!	+:�~8�S�'���r�v����]���S�j�[�^���x��IlP)�m��nC�,r���Z�]z�(62-��q�i���l����B�o��Z�;c�f�bU(N��5O�|���~�	efK�r�<斫�j�{7
?0���̤n	#K��MS���芪�F��|}->�o;t�V�nkݦ��l�;h���2�^!|��C����S���C�k�u�1G
M��>��ٺ�PW����7�W�%�ߪ�-�a
X���V��)pm%��O%��0�RCSv��6�M�u�?�-�^�hg�;����M]CL�66�t�7�yY!�*��
cw�^��|6p &���Hx�{Q��
�Ď�6�5
L�9X�:Z%�#��L���������:�G?K�������q�o{�
<��pq>lI�����? �c�Y�b�����h�<���-:�5��[�)lp_H�5?��@�Oh�1ft<%#�.��da��o�:�
E�	�ѡ�[d_�L��X�&�'��a��H����}�������N�0��ኔ|�%�eG���	��ufg7��S͸n��K6�E����c�>w��Z���]���'�k4v��r-��3��n��u�}�q���؃���e�(?����
�a�T�f2U	��V��,pL�9����7a
���2��Y�Ϸ����ge����r_�"%�ǧ���T�m�yN�ɘ�H^����� [��idA�}o6�����a'�9gI�ɆL�"�!9lԣ�ȖC`������>����^q��������h�_(�5�W �k(���,����L�7�������n9is�'`�|�/���! Jk�Ri�&3މ�6&L_�5�C���6���xt#��4���뉂��[�=��q�/��۞R!���F�$JE��%�-��"�Ƙo����fw������.�"���*�^��� |-��e�`�~/.�9� ��K�����7�vhP� �N�֮@e!ܚ_��W6J�~H�r��;����s����">��׊Eb/'w�^*�]Ay����!$(��vf�	���3�uD�3	�}@V]��89�!�2�4Ք�tgzݔ/���L�Vc��6�j`����"4����#���Q�d�X_ 7�r��DP����NG�n��C�"�u����i8����+,�ɩ@R��t^���@̱~�RI}�Pj���_t�G��{�#�s����
M2��/^�1a3�0៎����Υ���r�B����L��x&M�%[�?{CX�ͳ¡�Q/��P�3'����h����M`+ Yw��3���p���N���=!�M�*s]q���6�#�N.��"o���4�&���Az���GZʦ���a����k����)�%�<�Z�lq6I~`�m�i[&��Lq�vJ}lĝ�.��c�ػ.ςIU���a�ʿ%KaW�v�e�� ��ڵ��T�ϣ2�q�Ug�?p�|�y�Zg�72g�&�0�T��]�k�.m���OO F��A��e���b�f�,r_��t�ag�3_����kV�xY��I����F���>�I7B��z����,��uTt�_'%i����%�Z������4m�������`�Z�/�]�+��-��h��3L%�Z�K���������1�y��-�O�d&���ℑ��g�" ��+�,�ԑ[�{\�U��t4{+�ƣ5u�#G�����\`���K<l'�$�`����j�
��6�w�!�4����:�
�Cm���ڨ���D��%������u3�/�2�*�.(
'��3������>':���莹wK�x/
^���]�����8����7Wř$�9�oB`���^j����ǿ�u�x���w�~q _���Wt#�G�)�����0$r�8nq����b��vl���V�:������7K���ޓJ'f���Ż���J|��U�"�g�Pl��Z}R�l�����m~F��_:8�UF[��� �zF��������K��%���Ҡ'֩��>0g�t��5h*3���D���9�i1i���rC��]���t�ܶ�[W	}�KP�X��'%�Js�N;��_?+ ��*���%ׅ��nTed�qI��ȽE��\�_�-n,�4pGl{
Rq6*�|�f99a2�m�dKa�E~�G��!{bꖏ%�pt^E{����#bV��� =�\�v�;��V6a���sH-��3+7�W�^���x�P��%sB.m8]�vc=���_�:/Wf޿ؖS��!�����_>�n
 {�ֽw`��#��V���x6�����e��4��{\xmCB�i��1*�LU������y��W���G	PD8����f1��VY���k=c�ƌ�4���%�q�U0/�%�h�eK~�\>�M�/�s<<iQ[�Ѩ5��f�UU�v
0j�z5�ֲX ��4�@]�����~�$�����?HF��ԫ������k 1�ġ�#ᔈ�>���e��z9 �-��WB�/�Dt�)U֤>��uQ���*[/��!O(5H�tR����wi����K�S��<,�&�͕�}�=G�K�&��އb��txw	% Qb�`x��1@�P�K�x`�KH��_�4[�ӌ4A��K��U�r0�M&�	��{�:s�!5��(������r6�j�4M��ݘ�}�rt�{�d�-�~��� �Wk�7S�#�9?ԙ��F�%��b�h�r��w05֥��Y*]�<�k�w��t�ڠ�l�'����)�X���y$,����w�Ѳ��X�l ���P�Ȉ�M��a8�%���o������,��G�����꡸�P����'ֺ�I,��Ed�S�׆;O*Ʋa;�����������ZH;�q��7�V��S��nB9QǼ��6��u�K�H� ��lo�}Cp�����;VQm�z�� �`���~5�����I	^��V*i" �G9��OnO��i2�Qy��x<3�6�}�~��t��U�҃Hrڬ�$��ǌ�ڻ����'\��t�޳y���6x�L\�7�����nEu�����Pg8���T�V<��kT`��CsJ���Lucv�D��HD�L��΅oA�7³����LD4�>�#�����HB��V0�Ѻ�1�5����J�~C���Z��h�\��L��Dy)KXV�f�^���8�odA�b�4�����v�;%�6�j����x��?�9��N�^�ů��ʫw��Ì�%R;�l�v��I:'���_��4(�@LM����ISeeOyF��]@�%=#\`�������\$���7J��b�c_�0�w}��J�z�gh�j��Eo#Γ�popD ���N�ϭ�_S؞���̍g��`@!*��q%X�6Nn��J��f]:�κ�X����ښ�9�F觽���,�@��T�s[�av�[�O,4��6^�Bk0�K�8��[Zn<�"[�=8#������ja�59)��ao�a2�}<�)Tƒw!ho1���t�
��dK�69������t�,��*$��+��э"��>X4���j�f>5�\�ou����Yvz�v�	�~����w~YY#!�ȥ��L��VsZ�����c)��T';��4ຕ(�t� ~��*wy�Ccӛ���*Y��G2�{`f�r>�ٝ:h��)_ �(�[��7�t����Y]ԟz��w�l:���H���_p�7�2����^N��ߡy�u���(�?ޫ~SUd�7��E�<<��7��D!�t���Ǭ�f���gڴ�/�T��m�W��7.B���*�+kx��x.���H��f,U+��c����*�}���<k���1��%q6�Fc�;<7�����Q��U
�o�d7�����'z��*NN,J�:��
z�Gc8TL� +i�"y�Ю����v�t��~�8@,2����u��j*�$T�x?=���^P+Q�U��h/�d�P��n�h�˂������$;e�}���S�ٺ���q���T;M�� �Y���&]ŹnPXx����R&�]6���:�u#���<�1SVO�t���ݫ�Έ�J\t�)��K\�.IQ{�R\$�}w���	Yr��Q�9�>&�K��~�;�f[�F���g;��Koҵ�~��6͢���ħ�u���.��)w]�ch�n�x��4�z7�F�E��&�6�j2���%P���+3��~Y��I=ʀ�
�e���U�J�7���2+!��@�	'�
�Y���8�Ġb��z�������%�C5fǺ/����C���ɳʯ�����<O<�u�ٔSܟ���K�F��cv�w[y$�bJ��Y�m߹���B�DK	9��1���`��z�C���l��4�U�$� ��ύ�Ig��bF}�0�SF��as�Ex{&���-5 #W�e0�/`zP�O�|$�G	(��6y�a�2��@��!�V�VK�?��9�����6h,�>,�	%��2����H��8��~��ڃ��p�a�l"�|k��q~:��'��S�y�wx嚎�z�9~a�}�P�˺�I��'>���)�a-,��t��<J���US��>=v�1=w6sh��ܫХ���e�!���m��7�@=�j��<�X]p�{ ��Ifm���P��,�P��*����"3�?!Ep��+o�&q���7���`lA�[��8�k=�>�.*y$���*e~��gH������Cr\�و�aE��S.��|�[ES�&D�<���'jZ\��QZcj+C��[��T�u%�#���XkT�_b�Fl��!*`
m�ߴ�č�v�6�sǈ���;�
�_M�+7�#��P��{����H���l�hJ�*��\s<?��W�C@��Kvtv�@ɶR*5~��X$����3^G�a �i��_�&ι�m��nNw=ϪU����bS�����Q�² ��Vv�Ib�H�?���g���u�m�k@�fb8�$�.�A�"@����kEƎ�������:�k_�4?�o�����<�c�[<�4���W���(qs[��ى�2˜o�������m�פ6�PH��KUd�LH^���#�M�	���J>�SYE-�nr�*T=�+��W��l������
O+~E�`��q�D��0l�йw"����eZt��ëu����#�sfɭ��k)܀��\Z>�((�n�6F� _,��n��M�	V�6��g���s���R��qٗ��~�d�N~���N�2�N���{�Lg�C��@l?i���nP�������^�Au��]�(� �\\����ꁺְ�(u��VT�Y]�4&�6�O�~�SHݸ�!3>�ma�U�`'~6Lq�'ycQu���΍���v�����~5>����XY덊����_�����[d���G��b"�h��ջ�"�s �I���2@��r|�M�~�[���5~Y�����N��g H�8�V)������¬��e{�����Cڣje�9��,�O�����M���`
��ErA��v`'�:/�'fԾ��0�+��&n{R�j���̎��_D�<{�&1���1��^�;�{G�
2]�(c��߼ᆀ�2�K�ܕ����.��X�]���H 志�ř���3��a��� #y�@��7��#Qa�$��'�"���-o��F3�h�6�9p����L���!���d��P�]O�MCcI���50��t������������Щ���lV�Ri�Dw\f>-s\�x�	�0և�>�3�\�oTe2Ɠ����l(���������6�(�j�B*z��G�HH��W�A�����nc��Ē�*�@\!6�@�c.���l9?,�Q�w�����/��'�R�:B�3$9\����YU�6]M�'F�&妩�ʾ��~n�kϕU��Ƣ�Q���%_L��E�M[�	��h�n���}��t������8��fQ[Οv��$�U��\�t-�š�dcv�4��~�|�bG)!Am�4]�~�"�)sL[]�5 �	eI%�E��r墽�2$�MO�J1o���ێ	cX����C������v6�'�X؎�4��T�}�4���§t�f��\��������$pu7�	�hIa��4u��j���f5A�����[�6�8�C��*��upo�>u5�&�N�v������gQO^ͥA��"�5r!%��Kդ�v�����n�:�7#�=�nW�[������ڂ%�H�'���w&'$3\�s�S��@@b���h~˳FKQ��JV�*]�ڨD��	Oٝt�L���7�4y8�h�ζ��_��y�o8E>ɪ
����dw��I/�Æ�6�Y�r��#9(U�׋p�]#�� dשe%�I��(���cW3��"��iˤ%.˾԰D�C���s[r�K��ز]������o���z���
��?O�l��^G�9
^�����@f�{���J)��~�ūu7�w����a���3���e��(o_�j���͆�2O��1'K����YG���MSơ2�Q"��!�C'.=;R��/��� g(i���|"+�}s�X��v/�%��x�:-0ⴑ��kK!O�s���2�� �{���>��4�cK~1zis0t:
i�kĉ�M[�I�!��ӊae����M��0��x�}���?`ƒS���>��wN�7$Q�F�S������%i��-q�I�7�)�t=��4�
R2�#�P��[��b{w�������p�gtA�ACⱯ�O��M5�"P�GL)dՑV�SNwVRl]$��M5]4m3�{�����p c���4w1��I���̚ʎ9p�\�,��-д� C؝xOl��~o����a�=�A��V�PJ�D����("��4%h�9�g�{*�Tq�.y�M��p�����}����ߡ�s�dك$�>_���$�C5�r^�O��zӈ��fJ���H�嚜5�Z}�{��E��n�?#ݩ�0����<ݶ_�)��"{��5ع��e2|�fPl:��+�Ӕ4vX8��Mr'/�rq�"��Ө(��h[�'�<@ڶ���@�V���٤�>����-���"U$]d��7��>^�����u<�}�j��̑-`r4X�+	)S�%�d���rj�d��j�N����Ѩ�1�H���a�]����V��iO�cX�b�R]���A����g�_/��h%������I?\L�C�Y�ghKя�����6*!���v2vQ�R>�\]/����k�G|�[B��|��OLG��n:m���70�}5hQ*�W�VD�Z�D��o��^sK�S2H9��xXYQ=��Ӥ7�Ϥ��H����tڇ����/�"j�{(މ�@���r۾
�u�g]0�XDq�&��+�q(
/Asw��!��qMd&Ժ��l��`k�O|U�:�is��pp�F����ɢ)7� ���6F�h������v(#�g�+��!�#�dD���f`�
�Crn��*��U/�j�Zq?�s�(�Y�����r�N�>�'z]p��?�	Y���b4-�+�i�����c���y;��]����ϱ
��_�X�*K�+�i�5Dz��{�F�%�����
]D̃�!5�4}�����,��D�TS��	���
�^�-�7\�kK�s��w�9��g>:��zrr�O[�U��bO�D@��>�����v�t�(�N�UM�x��b�Ȗ�KX����H5=��]��k���]L�F.PC`�#?���π� �����}���X ����_�K����#��@,eP���!ѭ��X�%߮v�x;~���������_����)|3}h���6:'�����0���%�H/�dѠ��*�c}?!,HdJLir�dۂ9@����I3��)Ȅc/��z!� �;pzx#8"yH��2q�z��-���/�ߓ�0쵙��g��mt3D��7	yP�*�su2ߗl�����}��5,Rg-�<��5����'�Ec��,���	���Ŕ��Yxy	<8���]f��w:#��"_��m N&���O.�U0�*ԎI�_O�#�AJ�r�Ǹ���	۵w�U6�q|h����!R+7��Lu�+�ƭT,ز��h�Μ��f�6�q4u|>�G>��$�p�(�qe4S�䕈,��[�s�r.�%k(5M2�d���:X �t˘���5�s�:X�iZ&�����ݍAo m�0c�Uqȧ�c��ݰ@�M��� �a�l�d SH�X8r�~~3�j:�Y�w�`���@,��B��7@���)#�y����$�y=Ff�1�Ǫ-l/!L�w����a��~��6	�p0�Yн?�粋�E�ѻOH��Q�ݶpk�Kcm�E��ɀ2�)���J�CgƮ%�3:b�����[��LNc$\U��-�=�w��0��y�+�cJ,��#tGǸ���˾�|B8�n��GV7�էp
FM`wS\H�=�`�A|Џ%3��C�󽷗EG�\���¶n[gDt�<&�j�՞��Lz7H���{,䁪:��\��]L�TC�����|�N&&E+!;��/2���#N���?�	����-�2k�	6qt��rKv��Y��$�;��j*t��s�{�?����@�8I��^�Ipb�9��~(��;��^EL3-r��bߣ����	jwe���(�31G+Te����?�ktV`G���_�P�	3 �:��O9�5����u}�(Gb����<��I��ж�?���REԲ�F�n.RÊ7�z��D�ΘV�|�5�����:O'��z�Va�6�̦��!�P0bf������O�L;���f�_����n1��у��Q�Є����0 � ���}��'�**QO���S�����,�բ�w�H�OG�Αi��0��vợU���Gio�<�� ���ݞ�ѽQ¹[6ZG:�g��*�AUn��h�_�i�8��ͅN��eh��I�D}���C�b\��
P��7stK� -��Sl\hc�بW:l���A3)TC?�]L���fD�-TO8p�_sT"�G��T�/]�|,��7w\��#� CMܓa�6�6�K0�liF�x��q�P��&��.��6�������Kl���@� Tj�
lԄ*��E��M{����wl9��/�)�������,F�LY�c?_�fk-�(�1��jfN���#V&Vt��rC��Ƀ��΂]��L������'��v��5"0x\��#k-J�����[r��d��P��BD<��ڐ�cBx; <I�t�Il_�vNmݵ+#T�o�^^�f�Z���A��h5�2|���� ����H^[/7��^~fc�Y�X�m/f����w 
pO�B�"�fд�-�މd	��P��,	MЦ�o��mIK��eB���o�~<E��Dv�Az��;��փ��vQ[,��=��"@�4��ҳ����.�U���VU����"���B�c�t��3쁤0��!�3s���}��=�:�|���J�����-���uwv;Et�@g_L�)���h��~Dv�'�?��ҟ�F�)q;�W�̦G��t�����_W��C�B�8�%�)<m��oYCtB0�
~,m�qg����K��&�q�]�4M~��/�Z5��:��Uz�!���S~<�C%	��Y7i�p����oS�K�b,eS"c!��O����?r�Jܧ��,̀n�C��0vv�	 Wy�Y�ɻ�Q��RFr����ؐ�%�*�R�����*��L�-\$�ɉ���G�3��'���}.�dp�k��|���(G��#��_ٝ�Խ���L��,9"7�l�,�@��U�X#�k�/��_�B�7I��x��7Gc��\�_L�Q�(cr<wy���0��F�>OJ�PL�hJE}ࠊ���֎��z��@� ���� ��MK���y0r�<���(�%��4�>�R	Rv���Zh�V���i(�"��q@8�;��%��j��AY�ʠ[�!�u�'ڬ� �xoI[ ���Ђ��r�0�F8���'�G�)�hRD�L�o{��Ovō��.[�};�8G������V{tQ���-[��1��`��9���R$OG}逝IRR_�rـ@9��5�Nb��+�%�\��(v�"�����Z���{����%�cjZ~����|����	!�����A�FA7�ND3֧9�}�7>k����6g��^v�O�͑\Ѻ�\��a���A��9�{�����L���\�Y�;���Z��Wiyc�s�@)�p���VQ��oa ������f�Jamk'��~��K������N���i�Q���x����b��4����V�@���H*�S��ҫ���rr ���� �+�p��(�Of��������Y>����_s����<f����>t����j ?
35��w��j2����w<{�U'M8���2�96�_����y׿�4��G�Z3Bإ��tUI�[��� 06m��q^Y�MMk�%�rT�8�Ԝ\A������R�~��mrC�]�$`pG�g��ϔ��FXФ�����u�����+-��Ƨz������)���wV��Z?�2m>�Y	���c��{��xA�,�E]6�(�
y(:B4	��n�H�~	�@?x٫P4F�h貒6�VzTe*@��,A-ĀE�
�sޫ/)VQǫzY��[~?��U��y���+}�R��r�5դ;���N� eA�F8��kG� �L�ri�fչ1�e$Z��X�}]!#b����!�
9���7�ΈY�M��ݏ��+2ݎn=o9D��eΪ�̭��)��U�[Kp��hm�dH$����V�.;�PS�@qD�u%�v��������|^ ����)���ȝ9l��;� ݀�O:* �����2�m'�vY]_oS� �\�P+9֠r'����&���]��=W_]Rr-�/pw�����4��7���"����,
[�e�ɣ0�	5k�ɥ��I���xD�Od�����
��_����s��a��3�K�5���M�x.c�z�vP~H�K��K]�7 S�Y1̦%^�*��.��Ўƒ�'�@�ؔ�.N˒uOO��w^��R�����a�)�.�3cA��܃�
���P0Ry�ʢ�t��D�Vfo��R[CbD��F��\R�זx1��a���P$#�U��9%!�'��6^�����8_]y�����OK����jc����k�~���xA�۵����A��jL�Fޱ-�2����$)8,DY��W=���Vz/Ը���"Ι[� 9��Dd����&F� ���Ty�Aod.�~��Cv;��kX�z���"$Cz�7�'��ˀ�~��\�\CO׶^��5�S�t�,����"���E�����na����UF؃;�Yݟ�_�����p��'�mø�l���3���+Š��"HCo"���SO�(��Z&]*Z��J��sYK1b45J�Y�3���ٛ'�ƞd���cm���V��m���M3��k����^�n����c��ǘ��)ZU�Q�:�Fz\Ft��jK�xY���������*Xm��C�.R���|b��Voy͟5�Ę�J�v��\gs	��y;�EX��1?�-�a9 ���'{U��	�`�c!͡��@�z�m��kR�"�[�S�@8op �
�h
1�F(n�9|�пҽƶ�n�,B&����l\B��0�13,����V7
�;�#�Mќ���7l��U �w4��cTC��@0�A��������������`���-�1TP~iO�,���+L�$D�R]����Х�v"d;՛���������u:����>%�ia�T��F����XOV�y��ҳ���=�Ջ!�I�w�Z8�&�MȞY�F���<0�R�&78���p�`�Rԓ�o�J��Fhv :H��ӓ3W+*ox ��7s�踭KC�n��j��!5 %;'�P����~���rj�zH�5��ae ���$)���1���F���v�Z�`h����'��$�h7LA�t+�����\)Q2	ȃ���w�s�ܒs�b<F7T���l<�җ���P�q�w�!�X�9�>'�&��5���h����9{p�ʭ��^]C-��dvkCȔ��oF�NyM$���JE󑴪l�|���٤�ť���!h�?5�@O�F^�-G���]���?kB�,D�O�H�/=-x%E,�M��jB�^��(",���6*ڴ�!O���dl�\Q�}��ٌ�p�6�(:H���� #r� 	O��e��g���'�X�vG ȯ�mZ��!�YWB�x�tب�\&�}`�$������rÈx��-zeZ�%�!=V���@A�5o�4VBEM���Rk��4/���+��dp��e�������\�KϜ���l��إ*s�� �%���>���Q��	�qe�N��!厯_�#��ϸ-l�X�t��<Ի��E/Pc�Q어��3:���h���H�iQ�V�-x��-��*���xߧ9RM;�{ms,!-C�7G�|΋�Rz��un:�lv�*�}�M%��9`�N���)�>�d½wN7_��"�~��7��S8;~,�f<�S��`,Bn����5��(�`+!�N����޻�- 3��z<C��6������{n.�t��(���x!7܁}K�/8�vԬ�w�䴴�?\�/6��50{�|�9��!tU2��P{4|�H�
�v,]��}�c�,m�ej=��Ě;�;�,����<>1E�V�8:��T��t!��a�kF|�h|����H�ٸ�h��]�&1�J��2%�-en�/��Z�=����U�����S8��/r]�P����N�*��t�XI�x���cN��֥N���2%��Uieڼ�mǏ�t�vg+�k[_�e_%c��ShÃ)���	�=O�Z���0J?����Qk��V��(�C"��rj:��8��ǫ��)�Y��ߨp����iQ��5+{����oO�i�M�,]�S�3��}fEe>ٺ�77�kW����WU�-�G�,D�>Y��&�z��	%
����gn4���&q�x02!�|1X�������9W�~�{�HOokAI5�
SY
�z��$���-�v�JsC46ԧJ��OM_p�����>_�/�Ԯ߻��9��dv)�$'��3zG��5�|������M�4;�O�޺UgZ�~@�7���Te���֋�ʜ�JeP���$�/�׀|���//D��i!f�"�Q�4���]@O�rs�i�r����I�9�H1�Э_$�!���9/�}FqD�t��Eh�B���+�.�xۗ���Lc������~)�/�k�[^�C�Z+؃��{߻T��G�X+�S���$Un�ۇ��Vި4F�X�.����-]���%s���zB�#C�k�ab �\��!���Y�ґ��GFu��B��1sBu�:D���)��4Hq0СlTs{��J�!9C$�/8o�@t�
�m�Flb����
ÿ����\#� �"���nf]�5�j�l�a7�w��Q�&�� ܇ʝ�&�;kҬ�y�fe��!��/��m��$�Lcp����ؕ�=�v�'�i_`l��y%H�%�n��/q��������	��~L͸�xq����"�y�p4��3�:�/^h�p}�v�#G��u��*��6�ղi��/��Y�Fn������o������pGc�����%�#�
bq�'h�]�����"ѣ�=�0�{�{�{�{¦�H	��H�.���&2n�mi�M�i��It���~��n�)@�-(�z�|\�$VB%�J��N_W:?�	�L2ϋ�{�����fİ���\��J��Ɍ+"�~�ۅHW{Kp��A���m��lv�{����Ȗ��1�)������'=+�{�4����dd�^�Y�7��k�{���e��酖cuᱷ�P�ΪSʡ����{Ӷ<j�GD3Ԗ0��_5Qš�Ob��h�s#r�Q�w�6��g�ß�q�����b>�5��._��H�J�y�%��AN�N�.�v-ᷖ !�N	�	�t���`o%��M�#(�T7�=;���W[ME증���z��K��6�%��5���Y��:T@Dۤ���?9�c��)	�GS��v2���Sbʈ\�$|,7fY1��8{Nߢ ��y���a?�����oԎ�C#�J[c��"KF�_�g�+J����Ħ��ҿ
*b�j�m.B��;3��UB�@1F�+۟,�l�����4K�$")�r5v��
l��qp#Y9��=Y46�brU�ا�����~�w�S��P<��J�s=��t�8ς�[O$[�Ɔ*_�UW_��j5�4��/ ��%��%8�w�Ji� [ˏb"l�YNg��Y8_���z����ZQWx�8m�	 /��K��՗�+�/잖��N*�9�
v�P���X�@�tY{�jvf�
C��|`�pz���9
�".��0��P��J"F^��	vO�i�b�O_�t]�-��/;v|pb��u@���>b�m��M�8�����{�5�=�9ۅ+ĭ[�1^=��.<��XR1ߚ?��(1�?�(���%�5=�RXP�Q���4� ^
3�3/��ɀvd^�$���.'�_h+�l8dJ�@{7�A\0���i���0��×��UY��x�o�B�2m��:<�|�^v�"� l�K�p�F���ʔv���@N���m�ٟ-�Y_��m�5Z�>m&�>V�s�84����F��C�dA˻ܻ���n��/Lن����8Y�ܧ0"��3l
%�F�������#N_A�/�5`�v�0]!9�P��:����	���׎���"<�w�>9m�S�w��y�O����V� M�Ə1;#���Pu�U���)�V�-������v�%36�=,��~��;��9��&�'Sg+�?��P�5��Lܚ�s�)�?<�u�d�ߟ�ܭ�꽽uP(�X$3έo���(ߖ��@��%�W� izOXv��2�<e��匷�5\�[�O�߳�&ބ-��t_2{�V�FC���f���Ȣ��y2GG%4h�c^0n���!Ss�~UX�*B���"���Sg�� ��z�H�A�T>'|��A��ق��tƘ>:=X�r��e$�h�
���-u�f屬�F���7�K�5�c��Ά��'����=G���Uu�����+0�U�F9+͕���g�:��|�Y<��i�Ŏ!���*�4��7�\31�[��14�kz�s���ީ���Y6��X���PRLo��,B�^h��CN�y�eoZO�����J��v��I)(o�n�.��H�b�<<�:�����ʢn<k$@��
���\F���ڢ���W�qk��<��s��p����U/�
��H���lQط�_3O]�|{���f��㹊�������n:�e�c�ν��$Z���
T�ls'��_/A�Cn(��h(E�0V��o�q�5�g�dle4f�v���qI>,{.+X�?uvJ��������Z��T_��1=�%����W��Zr�k�X�n���������G_��Q[���|��ް:���[p���<~�j�p�q�]xzt��d�H�4�!A�u��l�L�J,��"�E�au*��
��lZ
qq@�X�����q��L�9�=����t^����i��B��M�v���,�MP<)���G]�Y�G?QJJ�?hl�c=��?"�|��AuYX�&b�.�� m�Q�Q��Sa�W���V�i�x139��Q��݆`�צ#If�su�X���y@97��B��ԮݤىտįTb\n$I.��'$���Z�82_��Ż1�	|?@���]��I�)k���DRą�cJ��U�\:�yǌz����r9�p��*m��X�	�(��-t����w�f�������R~hVj+��؊������j#ߟk�&�,r8%�8�(h?4�b'�0��yF�U�zk%������6	f��|L{=�it�^��{H�jԮ��}'W���c6C��]���y(ڤ�_~�R���%�	�(�!��7�U!�h��aqTwz�����Ux�'g*Zx)���X�Vh��g�"�� #Vv�')���;�{i�@����Ş(I�9�:�a�!�M�r>��Ȥ/*��*�GR�H_��L�����!!j䏠6/$�OY[��Z��y��+V��sP�.�>IN
���,��Ss$ZbU��^�&N�����%��A��H�.�⛡܂/L��!�ю5�|��Ӛ��u�+T��oV(�x�>t���2D���먐�C�&@��h`�޹�E3��@��[,��a��ľ���1�L�V���'��ikB�� �.��v����7a�)���b#~IDk�WK#�5ި(�]ְ�<���!��}�ΊoW:����[,�U?M�2ڋUYm�-n?ٙv>��q�Z�17����/J��!�hyH�N�t��Z����|O�R�����r3�]�v۴����cĲ� �Ĕ�lA�m�:3���4���P����ڦj�ܸ��-p�{��Ǿ㖇��7|��<�W�~�5�~.:� f!��r6�˱����k;�f�G}����3���K�����]'���0E�����,�xV����/4N�)�K̮�Y~WG��b��ɵ�s�Ց$��8�P��LUVe>�C_����!�f���u���f�@�)��!ٮ�`x3�����|���wI��7�*hJ�k�S��-1a��uY����':��ى�j������mfA�\��ZW��O��΀�ŵ����_ߚ��6 B)5����JTD�F��Oh���:T��	�[��rÀ����<1c
|�i҂3kL����/��Zna�ְ.ky`�ӕ�f]-r���mp�O�1�OMq�zt�"A��d�������䎌AjuUx��6t���|8��ԍFR��@�v�� �J�5��\1J�%� ����̞����c�p�fҪ�X��$Ty�p��<J�Cr0> ��F�?ڵ~���)$$ ��o��Sq	3Q']�R�y,bF]�q��[��^|0��?��,1���5	8w�WH�r��n�y���9#!(5w8J�NzBV���E��6@��>?�
�'7g������0�!�0d��՞~�P��H�.�W�ڴB��V���do�A��+����*!8�V�,__L�!��?�l��x݅X�9R����+�H��� X�*=?�6�%H���Ʊ̬�J���~��{��s`C�K<(z�_��|�}��J[�Xd�lM�)��ĸ�I~�)��Ϩ�b#�2u�F�p�;�b6�w�^.MM>S��Y#��߰ZD�|VM���uN��s;DQs4¼�N�@K���e����~�P#X�jo�|W7['k�zݣ�P1�咷pqǊ�L�\n7���(�|��1�/�Z��GzFp���v�gg���BK�Sӿ���7"��.��C�O�EbO'�p/�Ib��Q�eCI��k��U�d�V���p��ݰӧ���|E���x��F �����.�gj��u|�%�����SDk�=�z�ĳ�g�Z�<�2Q����ߘmH�&�O��^C/���i(5�duM�82+ONeY���4K�)����>�������3�5��� �� ��t�����{<�sMX7!�$d�+ג\�u��o;���31`9.��V=��*=�	�Cܳ,��]`0�x%�8=Ƣ$�<�Mt+��J�t����s,�`�l�R��B�9�����f��TX	y�D�T�rN:�3�MY����>4gƦx����פ�"-�K���{��k�
G� �TV�89���"��6^j[��H]d�X���Nj�d��B���t>��D����!
������Ή�����҂Wo̯�W��ރέ])�G��%������@�ph�#��be��VaLEB�(׃�	� Y�u�J,
����-�Ē����^�._kN<��0�o�Q\>�������W��69��ʈ�f���T_��v�XV���m�K_��g��S����s�N��F�$*l�5K偖��,'���]�1$���=�z�,94����*��H6W46�\X��>!���J-��r�ǻL�TG@�¡����d�,��ڮ��K����G�����V8�5S�v5�-VL�6���;�2u+%���=�zľ ǆ��]]tB��<�3f2��P^�M��7��U�sY Hz/B>��s����߱��(S`7���%���Q�?�ʹ�� �1h�A��ﲢd@�`)���0���7�*�8%\9�fY"�A��`;*�.Q@%*��p���e\^�t�췱P�l�UnR�D���[%���{������H���@
{9�Kv���W��a;ה���T�a���)�𢡊�</?�r��F��0*u��j��kDmM�^Zݕ&ۤ��}R�e-�`�>[���� qO6v�){���Fg�R\�K��|v�[K�,A��<��6�D�%�ܦ���j��u'�6�G8c1C�}bca����^ٞ⳿t��`�6U
�}[�s���O�i;�7��B,˒!J'�gX]�`PK|��\�(�;�$����XH4��K��>���;%�՘DB� %��I\¥�]���#h�'�uրp�G>�l;�v$�pC]>�hUE�:1+�����9�E_@������_���b"�L;��]�E�	���r�qǨ=���Kcl��vy��_��ͦ�E�<���69�)�DP)�NmgX9�o�{��̢��u����3�<��r��p��)��șA07���b7��vo>l�u��m�p%���+��ߺ�S�L�S�T��Z&��=�5s�z��a�����c@ri�0�ݦ`�,�:c"s�(iǺ����i�,'�v�@�a���(1ś	��$3=F(��CÚ?��f��bx���i��kY0P�aa�k2�d�gp�Q���`�pAjE˺5��~�u��.�!�؍&fA:[�g-^��*.�Q�H�ޜ�}/7��aPe�V�zG��}E-���B|ţt�9N��P��̙k�}�P޷���ĉ���Q�Z����ӽsW��5�_�'"^�Tv
n��c���eu���F-�ea8��j
ᅇ�8E����a�� �!d�*�-(��[L��T���` 6���:�k䋮��"l���7ɩN)��5Pt���6\�
�1�ȣ@2�qh�9w5:��L�8]i>������oӂ�y�c#�8�j`���C05���2@!*�^$R��(�k�%ZЪo�8�l0�<��_�ԐT�:���Oʺ"[��0Qȅ�T�)��i,�&'�4�CTm��i���Y7t���r��W3��@�'K��
��_�N\�!x�^�m�xͺ�p��ܴ5:y�S�?D��N��7������$��<W!�S���#��"p�F��d$�;a�Uc�9�à�sGh85���J���FNt�u��������Jq23�k)��W,[�{�>e�#�~⶿�,�7ɺ��9��J���s�����"��)�#�5_��%��O��Gd����%�g��a,���.UE���3�@pb�ؕr�3{�Q��ak$J)�i�0!�B\�(�:;"U^/q"|��V�k��c��.~�|%�FCJ�4m��}�J���پ>�q0P�y�c����"B �!�mTt��tb�����Y�/s>��a�&���ߢ/Ӳ���{{X_@D�=I�ޱ`_#)��D����3���XY���1�Ԛc�x�������}�(�����et�v�+vA2��w�OÚ���2~�k@7Ǻ��r�;��嵒���BV���M�E���L��Q�,�:�p~N�$七�s��Ɣ�1iF�~�9ɦ�#����w���0�ƶ�n���o|������VE��6��.r�?	]V���|i�H���,�g�RGl�F�+�'ߩ���?N�~^䃐h����-��
���3���üd=ÜF �(Oy���y���r��F_L4y���Q_��蓅��0M壃g.Exy�Ld��@�^l��K�Sx
�7ٞ�$���������W���a�{�T��3g� #��Y��&��-��%���i��)��uQA׊̯db9���i�C��"�'�����R��������[1�9�=)u����{<_Vl��zhD���;]��f�_^�����k½��}>���5�-7Osa\�A�1΍o֠r@\J��k��������^�R��qK�2�>���F�y���w~3k�	MMF���b��B�p7j5i&c1��]fmw�Ni^]@�u�l��F��#Zq��Pb��ݶi�ܤ,�S6�J�p��/���i� ��g9l [��p~Z���l�hڵ�^�J��S���w4��cv��:�E4���,��Y�Q�^cfx��O1k����+����|{��v���{�W��8�<A-���.^+ӽ���r0HY��8�@'K��K_�BC�.���N-E#H�x��=�ݩd#j`@��n�|��KG꿏�"��I;��P��n'��������Ñs��c'�ȗ��KQ:ih�ş�dl���(���m�%E@�{>�]�9��gM���?�0&�掶*o��$Գ�*�ɹ��[Q�l�cY�2&X��[K�Qk9�����O���W.Y��ɲ�/�v���� C��S7 3f�'o_��aS�|�/�z��9BE\=V�y�Ũ�aI�W/2�4&�s5z�����7����bp����;ѧA�#�斿l6<��-�E�)~��0jp�y���{�3&����`�,l�]�p�۴��Dչ4��?��Lk���$�������T��� �c�F�D&��n&�飮�HO�J]A۾�"�c9��nz��EW���/{r��7=�F�>��M�y�b�+8 :F���K}mFbB�tw�Lk,��[R�9҉���	��.[��WG#���%E}�
�f�ݟP�y�lV�I��G*h�NݿHI�RCA��=ȷ0��Θ�(H�P^���K���X�r>�DLM[š� (�N��:I���[��iB�����]w���ɖӀ���?� Tޟǘ�}T���Ɲ,�'�qdK�bNi���v��Y퇃o��2;yzҵ�����=����BC�3��2��\�H�I!p/��@Y�z���b��~�? �y�������-�z��~��nO��.��%�������������K��Cu�K�2�n�&hi�"�mثq>g2���>}���UM[-��R�(q�T�tJ��oU����0F=�(���hI% �h�[�Q��'��+6��V���X	�7�Z�:t�#׵��*f(Z^!|ǽ)b�X�-9V����"^T�AbH/�31B^�н�g˔	�j(bk�+����C�Mz	��(4�rd�Y���d
��K,�4gW^ �5-��)�������vV&�/��Ba��~�o1&�if�L��Z���F���"9����z�3����,��~�J �d]���C~�ġ��n�
�"�>���eC�(��W�(�a�Nр�%�^�P��(2�l����Zڑxot�}�)�*�ոh]g	澘�������&��^!0��^��66ZTj_D'i�yw~��ϵ�J�jbV��ǝ�����![F���=Vb� Y��$���EP����1����j_��?Xv�&����+4�(���$A͈�� ���Yd����|����y��@�e�u��^��<Z1j'��0���X���?���~��k�#�Gp�9�;�<�]ȞT7v(seY,nEp�w��~n8�sJvH�*���S�5n��9�����]�9g�&�ѣ�		l�61��y�7��<-b�/�#	�|81t��/B-���g3RT�C����P�7H6�D3U~�㦇�w�i�Y`iL@Ty�C���nA GO���R���Ѣ��0���>+��D�s�@,� 3�Bw�D��R��X�_�c)5+;�����J�T|q�T�Ӽ��zP0�GӨp�ő%/{U�4ڴ�'\;hΫZc�N�fsߥ�
��������eK0���VcD�>�L�c؜Y>K���I$JU���
�|nn�M�9��I�H���f���j^l\+؋Ġ�D�]�5ؔ�R4_o$����[��u���'��{B	i[Ĕ���@�J)GC]),���3W��K�3�njls9�9�~Pl�_A��jM��[ ~�+^W�
}�SaE����Κ��z������w����+4���<��vc�i��T�V�a��8�!�/�9�\#_	B:�$U����c�P����4@ +8���E�f(z
��̃��z��CeZ����R\ՓVqa�
�zB�1�����1\f����NQ{v
EY���N�E	ia6Xs;���������82�UX�o�[��L0	B'�;�1J@&�jO�:�f@�(�B<�ǵ�I2�+��a�f�&�rSNd������W�A��C�
�'.�k�ۃF>B���!�[����=q�e�* ��SSE7�T�ĐJ�a�����T��W����$vx����W������Z��rRǹ�Ѳ'��>��I3n����_do�mT��X�f�����k�mf�|x��h�0P�����(�ej�+HEy�wƎO٦^\�<Z�oan�	�s/�j�V�.y�6u__��3��"z<���:9�����|��2�Mk�('�Ұ��@��1-�۳�$�x����L Ų���37��C�Ԃ��3�|GX��Z�.�$�&��ݬ(���
3�'k��H�����6��O�I�ܔu,r+uׅ����C΅7��^XP�ZR1O����C�i�e ҳۆ"K��,1�Z��y�Ş�foOsz�ϧF�Q�C�m!h�<���A?���gs <�����e�Z�B�V�@Jl%�E��}��M��L�I*�
$���+���2f�8���t���������ʹ�x|��˾��P�(�N�)���c!��߯n�K�唐�'&��yȍ��9�����W�V0�pي�4C���Ɩ���|�_�ب>+��9ܲ��[;�SB��=�R*�&��4v�V��N����|�E v[<J
�ڤ��{mHa�ғ]	^@C��:/���T�����L�F��	4���ɍ��|�v�e�_Az�T��%w.My��F���o�SA��+���,������EZ
��SrY��k+�|ZrC��HQG]�Ҋ��-�f(cⱉ=���)Q��$�px�Oi��?��VC#h�;�~<�:���>w%"�݊Iv���$�I���0��Oo���ؠo
�4�!�i�lB��+W�iv��8�ɔtI<�2Q;��f��.���e���ģ"ȞH}�N胰e�<��].�`^�3����/�m���d��w������$� ZC�ve�Zr�ԧZ� ��b�OT��Q$Ε�fiD��� �k���%��m)���f>���̓�{�!���s.v��h�x8k#!��.o�>�FU�]pY���Ӕ��z��R �׊�]ʩ��r�8�ǀ?­GB�dJ!��$.��ʪJ-�P��V2Q�~��U�����ly�4v`�C3�U7��W66;C_�c��0�]�
�x��+(�������9-����OߵM�jڐ�[E���fR:\��t$L�Y��P�w�1?�ϗ;?t��Y��u�rQ=4ɤ49k	���z=�ܚ�ZS�(���6�$��������[�Rƅ��$�!�����2=����`K�4�&�N�W+��N��S�#��{��5���u���N�g���@�2�
/��q�����y�7W��r�̣��h��hv���w�3�F}N��S�:�VL�U��n�� ��ʦ��&�
��s�VU�%�ӆ��?��u��I�����}�ֿB�4�ޣ�,���r�h�^Z�<s�[]�P��mI溺]��dRC5��"�����mˈ��5@��o�ߚ�S`e^����H*���@��"��ܨw���n���R�Gm����h[̡a�^�[��@>y����>��`�y� �ߌ.��/��ɨXt������8�Y�X�%MX�4vp�������`��Q�I-���%��Ov�r-entO
��� s��t3Uf�+��.$�-�a�`=��z�I+�C�3DL��vW�s��v�V[�B��8�mIW���}��q��%v�$��t���?('e�
�F���Q�{�hN�)xWQ�ڢ���E�?;�:h?��%�1q��
qI<�W��g���#��r�t���-��4j*%,����"\٢�����]M����	mT����ys�?Eq^S��>/�X�2���P�y�L |T%ұ�%�M�P>���=c(�f5#�i�"1 ֗RZ���Iq�2T���!�u��x�0�
��e�dsACsU ZA�2p��Փg׵#�����*�M�?�B�	1 ��C(�|}�˒��zr"&����!E-]��{P���j�d�ZC�Y��^d�sF6B�'%_x��{J�U�z��_Jo��kΖw�Ɇ�|+7�5T�p�'�\iD,p�%�k�5_j�[��+�`%�}3�I�^��`�BzIg\��y���&�k�����]���i��PU��,٣.��HG�ϭ���8k8	���O� G�kF�������Ľð.�ϲG�;i̿FRpJ����PC�&��$�\׸P�m�h�0���Ғ�@��9�>($��_׭��d�admA(�ћ���DD9܈vie�}L���wT���,%{j���vS���SP�+rM��~�Zݒ�& * �4�y2���߆r���X�{-.��Efձi),���5��� eLq��^3�@�30!��<?y�½�)��6���u�͊a0������s��H��=�q���#h%��oӖ{�rR,N�YS=�W����-�閚�*�BG#&�-�~�F-�������#?�CE8��ǲ��>��?J�qؔ�_e��������n}���;t^�/{$�P폛����A��śK_�PfGb���@�l	=	�3B��ɦ�Dd�4*%�=�N�����2������?e�ǡ�D��xx୛�S�0k�L�╮3��6��'2~+�����d��LnA'	����Wi�I�'9�
M��Q�����#��n<�3�t4����|�)y��=��\��<�Pe|"��^��y�=�K](�%�m�R� ���]vU#I�!P6��-�ǽ�0�-�$��@�Ƭ���v�j�3��F��pY���ȿuQ�����vo�ly@uk�6��C����l5�zDHx�0��Q>���Qb0��~����2on��2�y�okq(��@�/����&TN��lJ��n��c�"̼�j���7�_f �����5A� u���!������i/SH�af��=�qIۗ���֤�o q�Hx.�u������QH-h����1���9���#צm2�e���&0;�Y̓]�S�s��S���ҵ;k�1�Vc���)�"��������,t�m#�,�L�ʞ�yy�|�w��z�P>�H-Q U��,��/S�2�s%Q��S�� i}��L�Ŧ�����06���W�A�#��g���j��5��� T��oR��=���D|ɍJhm|^(8�sė�yQ���X8qF�"�bɰ�4Ӈ2*z���4��E:3�S�'��1�b>���ϟ��j��ߊ���-|���ڌ���?AL&K�Y�D�#gL���e� �<��v���D�3ㅞS�A1���m���%Ŀ:P7}�.:�*|\��se~s��~���l�R�3�� �m��za��0� ct��|�	��͙9�jɓ�j8�|�I�J���ʵf�/Bt�p���eITCV�E���ªm�i�?���������m��M��]"���<�F�?��?���\׃B�ǖ�C�1��M�WL�W��I�+��J��)��WB�F�'ֳ*�'K΀��R�fR��(=��2�/0�TxGTQ彙Eqw���+�)5�K9j%+�Y%�Z�bJ�9��-�A��҈SV�RhlA]�E�U#���D�L��|]=澦��A���/�3�ik������i@�9t�""�h
�1|���m��*T�B�R�wk��_�9��E\J��p�7�<�&��*�ļֺ��J2��pA�T��Jn����	�SJ�'�~�hᛓp��'��-���߸l���*8)&=B�M�rӡ  ��>������k�B�+�'B�2��l4t�ڐ#+�m�C>{X�=&�j�p��+�ja�����ґ6i���`C],_�̚��#�$�����#�v|Wd�nIV�mhr8�idA��Į�Ћ���b��	.�!BZ<�]	$>k3��2���B㜪2��H5KZ�*�&�jP��-�>^tD	h�zK~� ���im-���0
��������wg�hՋ+j����Z�ɔ~nO~�,Ż�.'2�Q�R���F�	�`�˙���`|{���T�A���"��F�vF8����A$yF��	���C�᪳q~`�Ml�
w!G�$#��Y����6Z"M���t���;o�H<.&����@�i�,"Z;�ꤍ����gS5���{�f9�{����5U�v�O��rf�W�Ǡm6��@	�����ڊ�����H�B�*����g0cF��;���A����eJ �=�l�]M6��9?������j���kt$<MQK\7�����ټ���("�]�\�B뉆�3��H�|jG8� A[K�"�T#)�?�]�-jC0������Ku���
7g�,�a�h�UJ~�+��`L��<~W5%�
���W�&~�y�a��$���)������mQ];%<q�=v�����"1#p�[��v�����.KS�*���\2��C�[�NA�.^B���wy��$�|�JF�`dϡJT���B��1�Z0��%�ˏ�@=?�#>���icq{������1�A�� ��r�<���-�OaO�-�����gQ��f1��"�O�2�+�sd� �X��;����҄��>��P<��jg|~�u���M�)��d(F2�3��u��g�khL�v�N�����9���`��������.�l�z"E�F�7Z!c������D1��¸� G��\L�X���7�&�֍q"���n�Gz�ki_������u�����릝�_���bֺ�e�,-kF�9щ��l���&��J�n`�#���ܟe����A«�"/U	�S��Me@������7c�O�����i��S��I��Ń�Eې�gĈPM���7<����7��qX�?wz?Z�[��6�0����Ob���#�) ���Eh�~qC�'�p�ǽ.��Ӥ���V�YJ|{��`���6��-Wn��r\;��W�i�)�20��+� ��U�[ALS�ٖV/��.�L���DvK�q4�иY8�ra`������N�? �[,�$a9;�4�k�8��.0�-��)�Fmi��7��ꔐ���A�^���x� d~����kAűՇ�� �^�͔�i1�,���='�|�е	�"��@>��l�� ��@M�J�@����5~&n�U�m�h����6/h6���#�n�(��Ғ��3+��3pL�d����R�b������+*/���:9a�oB����{��v�l��y+�y�H��(���f��ռǊ�C�H1�Δ6�U/PY�tЭ-��VmPGB�y���H����^(�"��:[��9j�R7=a�x�Ki�uwoc���������-=;�Eǰ��������'�ƌ"kW��ڄ�M���"^�3��6>h]a�t�9��T�-������%"( �K��W[�t��U3\���mH�|gꍣh�F��*)B���2�I���~��en=����ψ��3B�_�#�qk�L�j�:z�g*GaDt�kٍ�t����pR�� 0톁<i�u�X�޽-G����wqv�w��׆��P$Z-�Ƹ�:lAż������1O]����?���2 ��!����AW��F�쒋]�d877���`_EI)�E��)-dlGH&~��'���(�v2��ބa��Z�(瘛.��P`��e�߉��v;	Q�s;�����og(�{�����vF����G���Y;��W��_m�M?|�����#���
�Cʤg)�[�'����-�Mvr�"���F}�j��k}+.s�N�@ �#hp�b�}t� ��s��Eq
�g��}VV��ʹL�M�N�������.�Dq v
���YV��"c�9�w�x�}pR0�퀓ĵp�x�"�r�1�8皛D������/l���U�$3t=/���3�ߑܐXQU��uwݷ�dE7[i�z=��0������/����]�0���Gkݑ2��Y���G��IW~2�������2��դL�,-��G�ev�K���gf�P�f4v���Q��'t�{z���OH��w���_X7!���M�%l���]������eU�`�j��d,T�q����B��XE
{wJC�QE�|vQ �f+  :Mlײ�@%�W�-[_���E�@�b}%V�)����FH�ݢ2�����s��g�JAث�>��%e��%?�T���{���L{�i���dj߿�ɳ+���N�]ʮS��lWhٕ��VJ�7ʁ�W�f�E�OL3��qʰ{�A5�������a\b�0�����k�De������ ��ۑ"ƀu�v|m����_�=H��m?@d�aH�$b�w��	�%x(N*����-���;Lb*�.n�b�柲Q=�IP�v�GET����X�ݑm���CO�GS	�r<�e�'e~�xue�����w��}\���Y�C�����7�t&�k�ï�{�-C�x!�I4c)�aQn&"/�c���o�yNB���8�wE���}�5˙<L v�˟*�X'E,�"W^;gX��HD�s���@�y$J�Da������?�r��A�%�{���uk\ye��}�9l��򴌉,5e���%�v��S�$��gPpwKg�7�#�0�zb�C+s	3�ѐ��b�ep�o�o�:����LP���G�hYf��SܦE����೽���� ��]P�<�j9 2�W&�}>��F��#�)�&t��S�tG��<s1�D��ݰ�"�h�ґ2�n"xr)�֑�;CQ�������7��`S�R*�"�46� #勘J�Z�8���0Sz9���154%9E	�����N�Q1�R�'5�J�M{oKc_�3�U�����4ή��%)~�3����e}l�������M�z�4?E��,BRz1q�dÌ�sg*����ߔ�+� �sF�<Zt��͸3Hֿ��� �~ �њ����_|M(�W(*���2r-�����5K��Lo֡)�igXL���6�)2t\��Ř��E������٫�t�`P[�%z5���+���|�G�JɾP<�'d��%RČM+�F�z���݋����8�b������_�6N�`��g��ԟ(�6P�8D�~q�ê�*U��p,��T�x�$�,����w��Je&itC�L/��%'���(-_�C�W븳q�y���7�-��v��CdE�_�R4��R�>8�ʟN7Bw�K+��	���űY,���JTA'��{ �^��"H��-�Z7cbv�z	 ǻ���D<^?CKs��	�$����r��lĠ�F��Ȫl�{���o�d�τ�6B�d�C�,�B$VO��<3t��C= B|Y�²`Z�7�w��G��}��;�G��q�$�����$S8�LE*J���wg!� ��n��M�p�ǧ����G�i�P�Ië�V���vA1u!�q��0�v�a��ls�^�~2a{j���YqA��-4V?����ԅ���
���N��v��S(2�GD�H&d����/5Q\v�)�{j�lP��
q�B-n�濃���ؒ�����cx��&�i�tj��U��i]n�h@x��	��u��w�K�>:F��"�e`b6�U�:)��8���w� W|#�ꄱAQ�μ�ݩ�H�~j
{�L{Q�1W�'�iؓؾ�R{,���?��/�KbkT�t?t4|4����	�j�.Y�����U(Q���ԇ�9�=r՛L�[̑99Cj�
��bG������T��up�x��]�%�Z��?�X�{�.����bT�3�>t��JЇ���x�מfP�3U��A�V�b���\�s7�B��'Vt�;��	���>PM&Dwmip5�"F�P]2����!ɮ�M��w��jb7�Dn�:��z�eP�9��K	�fhc����"��$�=7��o�or�t�f�R1ݕHahG�8mC6:����L�ͣe|G�m�D��݇�^؞K��)�[Nc�6R �uKF#8N��u�� ���N*?
�E5��@�)�C6�Ă�jI	;���!�|���B�b�F��;^��?�$�!=�H���w�j�&A�];��p�@�lJM�î�ht� ~�)2}��b��E�
�4s���!����
��.	+����S�x3AW��ʛ��	)8&���>kD�ֿ�\�Z��X#6�ZH�94��q0Է9�j|ܹ�`�X�M
ϽF.*��@��Dz�H4+��6j/�v�8Z���ˬaHr�7�R�|lBj-��D1e��Q���s �#��y�4�q�s�(�����q�X���}��r�t�D���[uVi. ;��x
,Z���<s}wv$��Ɉ'ӌ��,$��S6��Iw{�!k�n`b�������6W�A
�દcZ��[��ݞ�H'�6��`(��`�� <Ռ�����?I���o�B3���$بC����م,�{E>�z���רq_����d9����wIDM�f4�����F�KELoR�seNY(�C,�]�
Է�c�pC�8?�;��	F�0�z�і�$�7�c���omC}nRd����*����i�7?va[��%�j���N=c6a�^L��ך)�Q���4��WJb̌�k����D�������z2s��b��.�j��\Iz[�5�L	r�&� �v#M�PژE��SJ��=rB�Yy�B��~o`a8���@!���d����e)�u��lY�}?���f4xcqwB��"\1�X�m�����zN-�B��M�x��O���Ch� }�p��505:������k^�ž����|�n�+��vT�[Un�0,"H+�D���
*� =�'^t�bU�e�LAԳ���J�9.�dTs�3{�ʺ�,9��l�_��]�AT�~X�l�є�>ϸ8��q$��13����ޤ!Ly�v�yO������}~��+���9��Z�e�]*�Q&qb��6��y�T����U�l� ]��&��[i���!�wa�t�'IR�l�OvavX�J��|�9���xֆ�|2�G.��ˁ܊�#w��k�1�Xn!�u�0 ,�@�,����1���(d9�N5x�c}o�DZn�=�k�
��{�GetĔTR�4�Ŗo���N	"�[BF7'��vI6gک��6��Jqv*���kL����!.�ж:���s/k�m%�
��!�)�4�۽U�~�ʵC��-	T�W������Ѧ'dHE�-K�1M��n���2`\F�ʩ� Fp�ˍ/�Dte��S�w�@���>�<C.k��uQ�г��O��
��\��]4~K�f�?��ĳ2-5���U~Y�į�f�FP��V��)�1�R��p���Z�N%�+�Ly�v�3��N���$���A�D�X֚*��[� ),J�n2�F_�k���g~p�	��h��@�� ��	�lv-��;�v���^Ƿ_!�MN�+�+
F�,ֺ�uyT5m7d��ͤ�\OR$�<&�0�^l��,>^���k��7JV�{�3N_]��ӕ���5��Š��m���ŏ����֚������2V��E�'�=��4o�k-���Ǻ�v�����Sv��
�K,��t�����h[�����lm �K�m؄�k9�f�A%J�y���1�{����L�uWs;�vF$R]�A?����f�]G���oݸ�ɯ]'�ĬρJ5�E �w%���4�3�hz~��L����h.���o��[:�EHn_	k5�_��é��LZLF��1`�lTA?�����"(���}Z�4L��q���g��i�%����.�����n��KH�MeD.7E:��ր����)w��GmfH��F��./yi�w�>����v��80����v#���d����a���J��"�P���r�0�T�J���`�NS�̈�m.��bb�HZ��*�j�?�[!�x�LS��'dkJuyW�w��\z�b��HR
�{%���Z��,q����Cr�8�`#O�`i)��P�)�q�w�V6S8����O2w����G#z����M����^��"��^�+g�G".$���[�6d��!q6��s+�p�c���>�Ȗ�S�?�5���m�{�+C��`���+�[ �-B���{k�����	R�V����5j�����mJ��Ha��H����)�.����&��lQ��_?f�����A�RGY��w/��d�+X���Q�`�#6�5�d���E���T`��4��m�޸�S���c}�����c��uP��l�͡w�S�q{æU�skS-���,�Tr��)��I���8���T\��u�$&���= o�5�*d�ؑq���i�� .�C�@'� ӝ6꟒Z�یug�[��(Ң�����+?χ �|�/�7�
0������F,�4��/n�t?�|��܌�j*]N�A�����]$^6?G,As��S�M9��U9 �׏0zSe�`&UN�g��"�xWZxI�-~M>:�s0���^Dp�,~�JF��U`w}����[��-
�;�̷�)����h�/ɓ������#1݉e\E�SIf�a+Y�d<���G0%��lJB���0a��fq���}�ï�<�'̀�����f���J���bק�*=��R���d}ý���cż�&vB\F��d);��nR)ܼ�̢�1s7O
_�[?��� ��{P�+�܌!��������@+������p���hfY.�ʋI�rqJ?h�� W�R&�	����8?�mBq�_0#���ۮ�>�O���(a6VI-]j�M�ˁŦe��pn4�� 6K�������; ��I�q'�0��w7�����^YŲ�ɛ�������0 �^�[��s ��7���ND���B�!#�^�Č�ֈ%�W�C_���`+��r}�,�Os$�P�pj�r2�b�)
c��6 �����h拷+@���&9���8(n���`{���a�`H~�6�1�1�KD�A�k�|�.��q]X�l�:�V�3�a8����k�S��!w�o�>�^�b�Æ�H��Z��W���᫾������s`"Vz�]�M�lpd�{f���C
H噦��
�!�	3喱S|�z�U�1�V���&��o���p�Sr��� ���	Q�O�&/����?���Xp)�6�#�:Z�B��x�����}X�B/!Q����ķZBUԝt�T�{lj��G�;M�PJZ�N�m�S��x�m]���	�@ggEa��R�XJ����r�����5��E�/�˭�!��s-Ym>{�t�u@a�iNy�C���k��V'�����c��Mg9���N9C��#x�huO�L��+�W�������$Z��dd
��+h�5�|�Q�<�RX�H�h9B��a��h���a����񍴍��S]�������qw��H������64�ؾ"�
d�������L�K��Iر�#��&�'�:�2$�_b��{o�̩�8[�@K3�/ʒzc�!S�v+#�����Q����T�=x+ ��	���L�p�f���˗B+4Dk���ܧ	�}6���JK�_��9j�.sy�+�����i���ڊH�|lҗh=:����ƼXh��RU��z���F�.�+�W� ��[Y V�U�ȳ�T�^tc/��c���<��һ7�7�I�^��X����X�n%��/������h�B�|����7�a9ܦ�>��Pգ~��R�./�:=��Yr�&k8�C��V�	�.�/:��3h�H鸯?e!�@�&���:ij��SqvGn��h�G}����~^�tQ��c�I����5�O [��Φy�&��R�H�z+��"�nVl�5���J&��l��=V�o0ڮk4��Y�Q��jM��Rd�cr;��(�$�۾j�>��6��Ψ��=�/�J˺�A�d�����X��7]	d���9��ʜ�cv���U���?�/��z�V��(�P)������<x'o�}����N�to�ݛ����sl��Xߓj��������P^�M��	���jk����[��T�N2KQՊB�σ3�@\�uY#s�����۵?(B�}OdbPۥwd� �n��n�D���2+O-���`�2�v<�v�N�G���"�r;�~�
�� +'�tKR0~�*�n�d�����j�n��.��S�_m�]����~�`��2�u�R��&
���*b�e�j�j�d�������LQ�Ω��^�r1�����Z�C�� r���o�CT����}�1[�:����#�A����/���e����N�sf��9H'\{�*������c�a�l���>.RTy�����Xciv�/�!�l�����)���a��ރ{�Oo$�4��7|�k��%j��UD�S��{���y��mGx��>�exB}\������?Y��+�cI]E�C�a�T�u�h8e�P3B��q�<]0|T.��N�@D뢸�c�HL�<M\œH��8��?����NfxY_�^���ң����%ػ�w����5,<��U��Kܚ&k0�"�/�ۻ$�!滖���[a�T�zs|���31biRs3�ӞtՓF��|���-�!bz�"7�n����@@�|���r�N�_Y�xU�fSVo�24ڏ,E�pd���u�CX펯��Θ�	�;~��4�=����v�� Umy}4��Z�"h�d��j�BF����E[�s�ܨb$C�� MKm	[������}�gO(��Y��������+��Q��W�3��l��D� �E��r�<ī������/�m�}S���d�sZ�6֐��-&iOq�v7�ƜK�*����V����t�'y��l�S�x���-��W]�Ү��Gwu�x)��&1UVPk������#�5��./\�gb�锳�¦�A����4����zK����q�7��=]�.�;$�� >>�sx�O��;�D�MF>J�~AN%��l�qr׈�b��z�QL��;��&�c.3E�w\�a��B�}V�
G���;ݭCGc�}�����	����w�땼�ۍ����ّ�E�D��۸�u�n��X����n�}�.a3C�&������#ˣ{q��*x/Wk��}������zr4��Չ$�� ��~u45 �|�4�%��p�m��|�@4���4��f��݊jm���.%�^ ��`�=+]��!pd��N�tOo�$AZ曗��Zf�]e3��s�zgXzV����< �f�rD��'])\,�U���
��M�8;D��ʹ�+Y�K�i��ձ��W~#���?e7ߍ�I�Rw���b�Gp��8� ,9��A��Q��q����n�`���<�>������^f�oN�Q�n_���}:&h��Q����В�V Lt������ч��(�X��6I��?�1>0�K��6�������e��=��+W�.�R����x
oF;�Di�K�}zr��|7�^�y�>Q���S#��R0q��3ͭ~�O�U�}�b�A�"('E�io�+����2��DO��.��*�׶H��ow[v��u��>�=֋pfAˁ�/^��T;I�u=R��x_�%%;@���U4��������ݐ���T���y�J)��2+��������}�L�&���M��)cRB��=\P�^p�NB�9v5FiE5$�`)Iܶ7�M�C�|�6%1�oO�F�jB�M�cj�8}��S�{#䧬�٬�_�i4��o�����:n(�W��B���R��l��Q��7���/�.��;$Y�)���C����Q3r1��0A��9_�c���5��WQ$'�lXb,��������.��{����v6�y#%��:'B�A*�{Z�4�Кǯ��!����H���C�r�C�����7��Տ���`�G�J���u��"s�y���۞{�`
�'S��cϙ�}��M�\"]��!�@��ab����=Ҧ{3�|���Rb��q�.}��Q�J�m;��ǅ�9���u�6��Evl��݂V������a�:�+q��|^2���m���RbP���ު'����qS��C셷(Y���9�D'>��?2�e�D�AG��*�B�H�[^<�SB��6d��L=�����#;�}i�C*�*Ia����7�Gz*�q
������-b�c�*kߏd<^�<5����w	,�
J�|��EXGsh
�_���m}w�d,��r����?�㘈���s8�����G��Zz��r@�j<���o��YD^���Yԃ8�P���EW����=�X�����g����^+N���j]��t�0��2"f�Jz�<B<H��4-�^�����A�X������xX.x�1�8�XZ��?K{$��6��B۹�܊g�ܬ{��C��(��P���J��A$'`�)��Z���My��a4�N F�z�� �	9b��p�����{y:�L-��A�����z�OnD��;�Ω�9�>;��+�S���hut=�f_ǥ2C/���-�V�%@�I8�R���n��F2+R*�-�w���A��mj���!���X���`ǡҏ[�daT0#�i×�-��7�TKq�#�rh����D�~��~jb�?��RA�2-�I!գȖ��sI~طf�
���X���CQ����N�D�hG
lڝ��(��>�Y�t}�~0~+z��!kǴp2�&?�K�o�L|
V�m�WhkMs�o"�E��<� ����H�'��..7���9�2���>fKBC}m�	���'zf@��2k��X�9�ODM&h��2��C����kr�SYe�����OFhTe�'�p�ኩ`N�'��R��2,��i_�U{$�w#(-ɢ�`����F���@������d{���n��@��*�Q�h�qө��Ij)������F��I��">4`�]�*�W�ٯ�p����r��uT���K���<Ə*T$^��#� ���������ғZ�ֳ$m)��J��uiҼC"��Qs��C!}8�d�%ԟa�I�/�h������&��$s�
0��/�&����
�D��Y|����9�{�$X�m�I�<G��� ��W&�<��<�|�����9X7�Ndr2�g��zSW��W�̉՟�H�,Y�$�"\j�Gy����@s>���R�զ�o�dؿ�,�Ip�>@�N�X�A��ew�b��c�K����P���P��/��.d��� �O=��<�Mw`xѤ߭r�G�V��Q^�h��Md�[������A������Ny{��H�Q���{��U�P�D$��Hu��LIs���g�ϕ5ꌰ�]�Ǆ�ROTz����s��G�^� ���x��fA��i
h?��Dr���U���#K�Tk�kj�+�����T�u%�D&�u6��]�	/�s�s��{�]�����|6�*H��N�(��4�ώ�J�3�P4g�D�olڈ[�����k
�`�=�q�N7H�|��l�e@� ������������P�$P$��g�u*��K��Y���ʸ�.G�T���I��Y��{�M�n�Ov:�C��"+�e"�o����,��ˌ>3	.��X�y3�f��(�ξ#�X��O�*.�3� %fP�n����F�X΃=H�(���6�%z7w��������o�#O�Gک_ݾk=��C�us�ú��6c���N�R���S�����c4��d�fmbc���T��v�n�����?7@�B-@	��O�Uӭ�$w�LK�z�:��b�M��r4�P,}�x�x����.���{��uh܍�̞|��0��	����׋S*+@g�xT�A~.:�yά
�����D�^f��b��+
��OW/")�BC�����!,גX0A:�L�Ȑ�w��EL��9��=����"b'
�������МH����gI����^}S�2c������B�b�j�ڸ�<��C�
ލm5F:����ɬ�����F1�;��,���|��6P�F^�6�-�����MS��@��~��Z7iX�W��= 8N��[��&(j�-������[���#�x�*�v�����	kC���"l���i��m����	EW���g3Z���7���?KU+����j�/�� K�{�Ԍ姬��-I��@�<�*���or�73'����`�l�>���l����]�4$�ƒ,*R�]z���kmsl��rc8E�F�9�7�b�UK�Gs�����{A�44�`�ȑs/8���W�9��?�	��gֵ�%��V_qгd�ش����vqթؘQ�o�ss��[�����ۦ�j���Y��.��J��}t���K_��شj�D�P ���<����p�i�W�X:�����_�P��:�%��++o�J�Yq�O�_	�8�M4��DM�2ƹ<���K�꾗��G`� q�����N�X�m? ��+��[���	h\ѷ����R�������p���+�tŠ��xs�	�����JHt�-��o·�%���Z�����Ɩ{���Xl���0်�|	c�Q��j"�Þ��]IV��s��Lk�z�&w��P��I�S�I ��-W�G[���P���_z*G�Ee�n��+T�ø�6��|4);���� ~%��q��T��o�P�oށI'����t�}���/�l�ʐ��QA��ή�*��Wdg�3<� @в��s��qn�
$�o�gT��!"��u�=E��y�P�� H<v&p�Q�S�|.j��w�+`� ↸j��;���֟1�KiP������v�#]p�Tf/��S���#X�B����"H���tՖ��\��v%�G����$��7���XW�:�O��p�d C��	q�(��|`ϓ�<Q'�L!�BH�,��	�A�<���!��4��]n��H}[��~^𯌟�Z��P�vz��K	���B�55�9��X{�v=�fP����uƢ�a���=��k�� ��+Is�2o2r��M'rL	��|��
.��/W�b"#4\R�WvY���]�L��D7*rYK�� ��3���3v�1����B)��V�y{}�t=�kC�5�Iȴ���ţ��-�]��汞}�y�HP�|�d2�l�ח]ڌ����-act�Z�D�J߈�k]F'8�}@ɍ2����7f�~ҮWn�^��b��s���i� �7r'�ġX_H�I�.w���B1�L�O��A��,$&�V92Uδn:%K�Zw�e 7.��F	�s�ǻ��49�rg>���w9(�i)�$�,��1�0w0�j�z��3��� Hl��5��&���j(p��ﰈ}C=�;�S$ES;и�������`���d�*<9\�x�2�t���փ�nUƐN��_��V��O�+E�ާ�vD�ɞꈒ9dah�3���L#4�!Pd!�ć}��'�fȥ5�O�m�� �q��	��m%�t;���Bȧ�5�1ݍ���6�l�U�[oln���˓#55��!���e�*���?�6���X�aC�T+���Vc����{��g\G�-=�K����_��l���:Gh�P�@�A�k+�8^3��xU"�H:�xY[b�mc&�r���˂��t�������aC)��>��eg@e��*�A�+T>C� ��չ ���HWE���W��<��4��.��Ü�~��4|,��5�@PE-o���?�Y�,f���L�?d�xgV�x�*��{(T����}�8�D���5�G 5&E��(�H�RVeƼH���m�����'?C�
0��+���>:�Ķ R�l�H����rbUM�I�x��{���h9'x�R�|�o��8�O�x�� YD8�i�,6n�x��5�83(�N���}�r��pyJ0URSm���8?y�wS�X�ԥ�nA�Hڍ9�����i5F�mQ�cχ����&X�w
V��ö����A��I��"���뮽oW!0A0��91o閑�wE�&[ҡ>��/��DN���W�^���=���Y$���X���gW怈�!"�jY,�)���<rUz�`�ΖήF��L�P,�����BW�g��߈��ߥƶFp�� �1����vj��&�K~�\�哟RV���~*Y^Xi㽾�ͮ긾��N�G�fp#�$�6T՘��v+��Y4��z������/��Pn��m��5�˵d���l�	����t?&ʲ\u�7">������o[y�G��B�-�L��52Z#�zVL�:�@ISn�������m�E�M��S�����x�d��@ʚ�
���(0�y�O�R����A���E�*KT��t�HǠ��?``v8T�A>�=n]c��_/0Q�Iޤ�GII��F���l���,���'AO�՛/�� ��m��ϱ�0>��yD�	�,�7�m`�@����R��{>�S=�^�rKD��'<-���v���џC��Գ����Y�|��f鴁���y�;~]�U���C�/��4�J�9��6�$�����-P�L�xqlsV�	��Q=�HYd6��T�%:�N����W�'"�M�h
]�iBQ�ȿ����K33���q;�Ey���F��J���CB������/�N�Ǽ�5nFʵ�0z���L���.!;��f@|G&��o	o��L�]�+}�^8JQî~�����Eٻ�M���z[h�e���H�W;���ޅ������}H��b�����-��0���I���%�0��pp�2�-���x 0�{2q�8ĞQ��T�_�r�Er���5��f�+���v ��w��,�uD�3ҋ���	ռ�
����d���2,H�!8I�f۸2V��}?FxU"���� �G,OY�$62�y�V��lrpA@�t�
1/j_�_y*]��6@�SS[�]��,z��S(����$7����^�qp��툸m]���ۧqW�dGr���&w���k��z!׷}ǚo�}~Kv��%;���3�ņU���D1ج�\e��^!�����J3���A�.���~2��	5}~�m�rK���g�R�t�oZ����v���S&VEG���(��_ޅ8+杂��p����
�_:�X��h���0Xw��Β�en�a�^'���E�8���>�,���T�`��b
/�L"U�܉sR�t��$��('4���t��ȗ�6A�Zz=�Te�.N����Q�%NDO�J��60�QL��+w���R�g����N�}r�c�-h��=q��I^�u�(�8G�x�����$��O+l�7�"��0���H�މ���X��;�Y��P�J@��o�8�h9w;dQ#��<	����'��>��r8lK��M��B��ií�������t���p��p�TKhT���ۈ9k�_� 0�\�1�R��5�7-4�K�X��K�3��13�T�(����� ��;*Cq�}BV"9���D#*�^��)�LI��L[GF0�Ԁ8^�(��o���1���������
A���R]02�x��>F��#b�����w������0�e�G�L;�(�!b�}��^|�E����5�xd-4���/�7�έ�r�u[���~ �[�7�K��e%����\)�p��+S����RC?��˸)oW��o��wG�OIGya��@�k~�f����_<?��e�7�i�z�l�A���s�GEa59������ޜ������MH=��O\u(1HvI�!��Ȇ�4j��uS��zX�b�i�/Y�_͞' ��. �DHۈ�'A�+d���%����ؐ��B�V���c���"Q@Oa��	NY)����Hg"���<��[���^X�������a �\��j`N.�##	渊���2^6�7𺬶��P�W
��/���!g����Ͽ.00��K��g2�(�p����O���mu���$��5�.'*����qmWBv�Ż�Y��t�Q";Nm�V1��k)���՛^a�R���<��N�z�p�c��w�_�b.��8�*m�Ǟ)�0j�d��Fɐ_��l?�}��VʤXj�7)�Q�4�3l�"�{�k7���j[_�!-ZN�H��ci�4�@$ɋ4�8��-�
�d0����=,��7��yL%A���'�t�R2��"�~����3�D۫Ys�@XI�,����\��Yy�
�ʚ��n���ShO��-lr�I��~>�s�+蜂�L�]J����L��Q<�C�"S��1�Mˍ�6sH���B�K�go9s����	���D��>��@WQ�u��2���q��(�"�ڤXM�3+RIAv�(�P�� jD"B��5�����f��Q;�y:�[���]R��Bht�{eBf�ٮ�=R��%D�c`&w�lq�]�_2�@'�sj��o����iK_�l�>2��+8p�N�B=$��{9z�v4[~���{�6�58QΝ7N���{`V��i*�At�t�S�s�����ɝ��+c��"��/���y�ѼDD���J �g0�uc��y8��2��4�R濬0�F"�	��L'�]7���[e�?T̃w2'�*�,�:�VD�=�]ӇP vpR��#���MY�i�=y�n	��R�?�HӼ���t2#5b�cB=���T,Q���i31�{A�_wI!�hǐ���O��nǊ�n�n�2��O����k���b1۝�q�m�ٟt��T��q�����u{��Bo�.�1����h���*�|!��%����ܑ�c����aX���R>�������Cv�F�6�7�F1H䩭;n)X}�gA���T	���L�E���֒�HT�Ugs��C ����t�&T��-X)ќ�)
��`·gq��S+�x�ps%"����h��d��k�6�v�r�md-���p��Pl�u�~��!z���v�@���,UI¡caI�氈�^��bB���{$rj���ɭ1�m�/(���3Yi;��ǉm��XV��nR�CU,��P*���Rߩ�{�.H��t�o�"�@�10�����9��$�.���J<ǐ �\�9>d�-ֹ�#�rC|x1�����̌-r��z��Q��h���e�X��ĉ@�fVm\�����JBhu`�A�)B����ÚkɱG1�M���ɬ���:d�ѹ~gwЅ�Գ7��73�:i�_�"��Y{�p1��T�Xg�|:���� ��1���S�*!�yɥ��1�(�t�7 R����,�G��1A�D�@�77Ui:����v��6�M�>�a���������@7� �D����א*V�t�ۉa�r�@hZ3P����y\��9�i٩O=>�p[���][S)}F�%|_�%���(>��HiFn�p��ƺgib���z��I�`����Yi���C�g���T	������kk�_�.���g�H�-��,Ѭș�!�+t�s�\���/��G�Ȋ��̇m�h��T��_���X;�"�E1��X��2�S�=�h�����&wnjz%�8,k�z�h��`~PT���-�M��GX��>�W�r��]�Y�|�B�b���R݌g�\Ңo��)ْO(��J*�O�A�m�l*�@�����.��T�0H\�Y��P�>�xN�3�^�P>���E�`���C; ��!��*S��!�?M�QË{P ˧��.��㺔^���l#ܰ��Z(�c�x��ڊo���$��OQ�xY���ɋ�԰1��kr?����4#d*�淋W1.#�	���S��
kQ������Ǎ���,WԆqy�W�2{�H��p�o�#�(���e#˦��~�'o��ek޸$���Xǰ&9^O�w9�L���Ff����n��<Ԟ���tO���=����e��v~���
�Qt� q�D�h��㤢|�)����{�U��Pe��iK�sS]Hf���H��;�1ŏ��O���b�s����6�p����}��G>�z�����m@?	����4�q�MԦ����*�g=!����ix�V��D�f;�l�i� Y��:?MrC�?�zJʰ�*�-O#��#I�%��I�*�3d<�Ԗq�VC��V�@��퉢|`�0�_r��7����Q=��.�\ńiEB���Jo��d^Z{�5���������{��t�^s�9;��*ys�\�{��R�H�:��q{�I����n~�0\$<��_�?��@������ܰ70\�Vq�� ��DT�`�iXQ��iQ&T�Ĵ1�K8���b^OH�a�z�\O���1�띑/�)tLky��4�������U��8i�:��g���u]8� x#11x���\T�w�!^dL,�O����a4��u}��p�V @Dw�l�?�cSG�p:���\�\���4h;��x�{Y�^@���B�l��/����d���^K��Ÿh~T� ��y�
,ѭ�r���k{?��v�=o �6�nd��֘9Hg��ԒA�Q*m�	�,�_WQ��ʼ_�=�@�t�D]�9��=/��; ������l��A���n���G�0�����]UĐ�P����3��@�ƨ� ?����́�E��Z��1�F�:��ޮ��(�qHk��J��<���K�,���t7�\:��ip#���t����ѧ:7,�;C,Q+�UT�Į�7�L���p�N\��-}���j��p��ݗ�aEu{'F�#�=T�*����8;��/ly]�;���Z˦G���Eӥ���/;�1/%1���<n�<g䧩�Zs��ܬjb)*�S����{LZ:�N�cϕ��F*�玼揽�B,�vM>T�#��; py�1�w+6q
V��~i�Rl�^u=!��2���&�_�Hh�?}/<���>v��t`�Nn����B^Δ�2!������r��)�('{+�������p�Q���K��h%���biU���-ԟw��:�h�r,w�A]���r��)+��[;���7S��u5��k��c�һ��[,9h�%���[�F��[�k]`��V��XGK��-5������.����Y��H�%�:j`%_u!��Ix˒X�p9�{�����J 9A�`:LԗT� I��s������D,
��us�F�J�Rԑ�����l1V�Haik�P]dh��׈r�^�%k�$�%ruD ����'	/���-7L��]D9o���Qq2�Y�xj����I����j����ͅCE�m1k-�����ug��j:���B�_��KD�1��51z�P鬿_?���)�&0LuOjX"\C�U�1$��.o�E9|\�>}�B�����ōX�z~L~UJ�:b��;����Y�6�0�*�9{� ��.��!�ޒ02��+���)W��+Q�����0%�eL�_�ņ9
nv@m�����&�玙�1�Ϩ&���*2��^��a�g�udʛfI��M�t���;J�WЂ�u��Q�
{9�O�!o��|tD�ȧ��ɋ\�}��M���i,<Q�pq>.��t�rv����Eu�22�L�tƭk��xIPx��/���aު�L��\��zjwm��^1���
'T!w	a<ۚ�U�k���[�����������,���ۿ��	G�t��g��:��Ѓ
?���w�S��Wڝ�+SP��K,��_��"��zɺ4[62�u�B����P �{��*�e$gG����8kK
��c.�v���ޛ��^?�,�t9�_Bz��&&�a��b<L���c�����o��^��z6\�������G�5�mM���rd�7�t�&�M�U�s����TRtX��ī)�}�[NC�l�n���`��\��}ZQk�c�V�!�љ[�Ǧ�v�.S�T��L�T�<���мO����#[L\M�|ٜ���(y�Q�
�6�	Iɉ�,���c�z��A�Fk��B�����Ne��8]>��|Y��C�������"�o����o�]�@TX��坂D�����)��DD%���	a��<�i�^PU7�t�X�k���+b.���A&ᔰa�b�|i�=�S+��I�X�q�������A�iv`�7}y�F!@�丼��9�!J���С��=���!RM�=H<ڡS�s��9�<����\�/x�W� ���Q�� 㽫�����R��e�|��ã�������.����p�J��jO����S��D�-O+��kf��c�l;� ����[��.�I�U1䱁L��$6%�ӧ������9��:����\�چ��qJX��J2�Fy:;�W߫���,�j�A�BKC�b�^�~}J�jX�C��>�H^�b����M�6�޺�UvR��Z������/�C�yH�.2#3U��r����M^�@��18��^!Ma��F�����Y��F��(O�{̆�h��������^T���۞<IL���e�:�
�4z������܋���64��_{����F� ��b��\[3SP��ʝ+��	ɋn��A�$ɜ�"�"��7Cy4�ѡԿ7`郪����t�j��Y Ϣ�h�U�I��v&+�k5�RK���b�3K�E �?�����i$��ަ�o��(�(>�[�`Tw�(fLd{�	5"n� ̋}�W
FT1���\�7�6�ɰW�T��9�8Cs����"�y��,G�;�
�	/OƢ�0tq*��y��`��ٱ֕���jl)��m�f� �?bǜ��t:n�i9��^+|%-S���a�'�����g�#����A��Ԟrl%�$�$�{}��s��OO��S�ѷ�oh�Yf�.&SD�/��c�Q	Ɵ"�ݓ.�B��g؅���9�fDbɮ�� [N&F�#wW��n�et,���m-�5l_ݪԣK���i��t�����bg��>V��p��6�u�rg�u��9`Y��?ҕD���.	���듼x%N�DM��唗�����G��� 
_@9�����P<�d����^,�tr�}oP����j)0(sl�)8�?�@L�� F�l4�K�W�����t����g9�huL���#l�k�.;T׬��4E2"N�1m�	���a��җ6����»��I�u����?�2�z*�F�f���S�O�+zE��3�8�'����pP��ϐe73]�.�2��2�:EF�nc�OEG�@��0:����-�םG���Ƴ9㼅���I�2;(�|"�Z�b�}�u���>J��t b-v(j��F:�J_�)��v�3I���o���u��@�滽=��E6�Y}I�7B)�6�W��HAo�0���o+J�l#���c���C�2g��V�s�c���F���ԳR��9�(K�Ϊ�ً�*����$;��/����Wq]~�?��.j�6��;5Z�� c��F�{�����)��A��: ��'���t�ݮL~nl6��l��9��#����V=o��1�U��?��H����9.��Al�^��;�9�έ�>gJ�( ľ��;���ڔ��P/L}�XQ[�ν5�{Ե����l�b�q�Ġ=5�I�x̬�l�&�SG�=>�Ŕ���v9;έ�
E���Q[��g�o]���I�Ԝa-1�vB�����- �B�8q�kf@fA�+����I,��=���=�_䍂��|A�7}�� ^�gPp�|��h�0�3���u��6��.����d�G5UN���X��l�NP����6y7���� _�F�iX'؃��吴S/FI�m���s�	Q=\�pw�9�(��E��}��&O@��{ĩ�Nd��Gl�ٿe��2���A�����X=v�C>�H�]�U���.m7;���IAI��ᠯv����������\.B���1IG^��Uz�ݬ�2��,�iC�\�ם|�`d�.L#��K��*L�b�{�IR���WM�[��ͳ��9_���5%�{q�NDA˭f�F�m֣dW;��dg�?�0^�QzF������}�q��^�ܺ���:`q���9�V��'��똤�<ݘz�_D|��E��M7��U
�����x����~�?a��]��Z�Ui-">�(R���L�:-�kg�ո�C���
)�-๾;��5�p�?�Z�ͅJ@��un����I&�tk���[pͼ'-�ݐ�_�B�>aD#Ȱ�=�2We���kcCk-�ߡS��Z�c<�A`ӿ`�%+*���!���Z���P�?2�,�g�Օ�z8�ܴ��3�*B�Ee�GDʭgU�ӂ���^�k�K�0;y���/<��s���s/�����.�,D�\�BJ@`)3�U��8ƴ�7��� �C�2��*�����Cu�$�!=w� �������3��~���e�_�|���5����&�n~B���T�<�g�&�o��r2�o:����}D׆)�|7�x�_:b������>�Ă<��τlW������b@;�y��BQ�@e��?��f�����0Z��+�);�d�&�t��(y�Wmg�A�1�<�tx��b���Ɨ>hk>�����j��ߓK�Wնr�v�ƿ�̊"3& ��H�d�w��߰s���渜v�J�E�����d��U3���0�Xw�|��h�i/	F�1�+F�-o�S��_����a$-9�x�˚�[���0��>Z2b۽c��j���c�w�:��dM��<� N�crhH�`�[���e{��KK�vj�j�o�j$NY�C��*��9�F6��(^a��&t��5���8{v<^��N�@>Dd	��a�q؋�'�pJ�|�uP�o2īn�8pB�gV�J;��DY);+u�r8yԭ��h(���Y�b� \*C����l�&z��nfx��[#ơa`�=D}Zo͈���/B���Uv
�������
�a�iJ�����i����߭�Q��f61fj���@LV��Ṽ	�h=����g�E��ԩM�!����	2��a��&3�@��T�����UR���痶!��n��MuC��T��ܛ�y���na�t��P��:��h��'�+�D�E������glr}� J��O���w�@	NA!ܞ@��s�]w�	�&�ԻO��;��:|_Z�N1�eXuW���{��X���ҏ/�y���5<{a-p~ݿsJ��,e� !����ZB��-q����~N�AC"�TD����Ztw���Pm��l�9�A(X����������6
(D�IO����%H�JÏ��*%��s�׌�%uugMh}<��8�ɭ;6j�giO�$p�QRQ"(�z��(q��� �9O�^��L�����;1J6�3�F���j��@�b�v� �uei��y	/{S�>Ȓ�o�f7��=~����y�}Ol.d�1���ȹ��68��t�
.)�M�`�3�Z�@��k�l��>߭� 2?��"�Aa6�RQ�:i#'��5f?4���Ǆ 0� N7ǘ�ǘQG��ey,��w4��<���Nأ1���Q� �>&�U�BVv��	܎�y�6LwhJ,h�g}2�Ԉ���F�o��6��<��q�f�聲��O����g@2�ڃ�\��fέ�%�+�I(k���e���^�ή���v>�+�l��=�����s�>�8��s*����3�'΢�u��DjLS'i$8ؙ�0�f�Eਖ਼]ٗ��<�]-$�r�uʧۼs?;�,�3$��FJ�z���#�,��y�l��M�0�)�6��_R|4?�\��o�_˅�{_AM `����KH��#֬��t�ʛ@����uy�KǶGr�cn6%�ț��������8|X�C+6����]��Y�T���0F��z��%2��X]{����T��R��{�2�zn��=84��J�T�05��ӧ�.�L/���o��{�\N�2�K��?y��\:�6|h��)�3㻅2�������K�5[�τ�[>	W}⺧��b)��}��s�n).o/�+_Z��8�S,`և�&���'2_5�;�ڬq8b��5�ԉ?�U��
�D S�MN	Y�Kr�3!�T�1���;����j'�3�!�[��\0E��k����i�Z2�=Hf���:��c�w|��7_�?��k^�xэ��y�7��sA��~{��E��&�qE�gBwu�4P��/�l[t	7�5�O�Pњ�`�{�0�{��a���Ϭ�����z2�f���ɍ6�rtF��,�|'�4��l^jG�1bfgs���V;����g��ľ	����j�:����:�Ԏ����7�YjE�-�맋�������z��x�D*�Pw�Kct{�F�������0�����ak�J)2҆5�ρ�Q� ji�'e�i���}5�QX��0!�����6��\�yl ���BD�(LX`��/�Į���~v-i%��g�R	�&�X)ė�ve#�J��Jȕ4 ڂ��&M,l˜��|3Í�/W��.�K��h���`�Cds�$�d3����_X�.7��H�2�~l����0�`����E�N���}�1���{/�'�e���n�}�:QTS�Ua=R�
~��F'��f˞�;?���(r��S1g��6Q�I8�ƅ$�A�/�F%�beFCֹ�D�J$S_e��S=�Tt�xuם�L�]FM�+:��s�P+�09�@�Q[���s�}����q��z0*ke2��ϫ���MqAZ� }�R����gJ����Db��Kґy.�Q$)5n�x���T�*m1W��0�! �dQ���,�>r��bN��5�&2.?�{���b�W�i]� J;����Q �؏��'������Kd��~7�
9U����#q��*%�E��z�r5�����%�@0�l̼Z�3,��E�C=kB�� ᵻ}4%k�c����M;� �bϟ4�p�T�Ϝ���pZ<Sd*�E>�4��6��:a�ʙ��Z�H;l�ߞ�(�/Sv��A����#X��% AM2g��t7tT�#�.�0����eR�^eV�̥���&X�_h��Yǈ�V��r�4�Եd��3_�3h��F��4|b�[ό�s��G�:��o&F�����M��M�lي�$ğr�����YA딁(h���4�����-����U�B���;09��ay��w;��g� =j)��OP\��U���c�bj��"��<g�]�O������6�${y+|b��X�Ӧ��	���D�vqi�����ٝ�S}�Mr.Sor���k.p��T�;� m��5g�Ku;w��`��蔾+�K6�;T���@R�ѻ$�/Q[��T��Zx��j�C�n��}�w����y�udN�B'A[a+�c�����ݠ��g [�9� �!��cP|�ȶ����F��ذW_�6<��@�ܙ&Ɓy���|�D�Vf@�sa�Q�K�o�+"�� "e6��������S�!��,����.9)���A������ϳ���l�(bOc�"�%g�!}0#%_�S�!0���	{Pi7��籇�[�a�K��J���X�rh+�ы�7hvl\W����Y���3�����g4��*��9�y^�' jR�g{H�p��I�H1'r(g����`�����#�2<����|�e��pk��Wb�Sx�G��
���K����x�qD2f���)'��셦3	�Iך��P���Y~	��Xv`Pd��k��4p��˽�b(5ۚ�[���tzx�}���;79����J�@������jo�tTܶ��/c!#���[k��U���τ#ԑjd/�e�3�ܓp쬜\�k��sc���#���#an��}�i��P�b����cU�=p<��˅���e���2=8�-<�>��7��#+&�c���(!�5�睾~��݊��)�h 0�.�]r|�9�&We[์�1��(۩}�,(���V�R� ���,(�x��~*�	�`&��a��I��6�v��5��3oͭ�����1�@}eMs��՛��H�!! ��/`���h�t%� j�[�7�2�RdH�0��y4S%�x'#_^LM_gc�v>�K��,��}��DʩI���_s�pS��1��^� gg(�����2�˷1���6=���#Tq� ���R�9_�5�E�D��X�I�o�|C1w��X͋����#�"��G� ��eQ����>R�z��s#ۆ��GA�����$��2�}�5�w�1�/t���^���41����|���ج������M�+~hFu�aR:ց(��g�cZ;�IH4��%U�]{;�����z�Ό6|��V��#�mR���H±�՟�L�Gh�\2M�Ɔ7�� E�VO�ᔴ��z.q7��&�a��0�����ܐVO>S[a>�"�N����cJ��+�Cy�v�w�{i����M`
�"t����k�OOBŬւ#yvJ �����R�ѱR��q4�o��)��5e�z��'���`�̏� ����nK#SZyR��6E3��y`4����O�<B�y�wٛq������ �#�6�MG��Ѿ��bvY����yӕNJw���Ù��_�Kk�

�Lpؽ����:rc
����g�5L�}{w:�N�H����'Y�k��Ԏ&/nT��0M�/����Q����S�2�{�k1;���g�Kۋn{bI��j��?T�P�'�:p�=���p��<Gm��!HDo��K��I������ں�T�%�pP�K��Gb-���e�)�K��OŤ����Ay+�� "�d���'�\IR�k���ڪ�u7A�@�*̹9���^A����TJ_4 �4ʑ��흘r'����FD��ٶ��Z�`�����R`L��C��(\��.����Oe,�w�t�z�}��55��?���������� E���VM��[�UA��:���9�n+EB��>~���F����` *���f�`�%l����z�<>�Jj��5wuxv��@��I{�h��2@�1����[�z����vI&9A���O9�m)��$2���Z@��%�k��� �˽�3c��̯�v���;[��Or3�Fއ�c����iTUW�R�^ǿ5I�|�}�[}4�*���Plk#�_�x�(� K_�x��p���Y/WŚ{	���H�Z��n�(��Ujk�f�L��=�3�h��W��!3/�C7t�n����od�����,�A���%8�\m�$CCK)�E�6�DC����ݎO��I�K>]��|�CO�=�z�d�[J#R��4["�A9�L�BܔHlôe>¯�= B�.���7Z�$L�𼸡��`�q�e��Ӵ�ZM�
��&#���'"&�&�Ͷ�#��̸B��k������.(1�44i����3hsBs�i�8 �J�g�r�\׋&
��0�f~iMJ��}�K�m��B����8M�|}�5z�=�ks8�
��ƌ`"�$3����*˃��1kR��<�T�#�x{T��9�ǀZ���u#�q���)w���j,i�'�$�~ؘ2I�{s�P����I�~Lf&UI��K�-l熕�$�-]�-i���2t��-�?q�q��G��W�c$�b��*��ߔN�!X4���%���89�A�:�ex�P��܏��>��uT���̓��8�SޏWОӯ��	p���	���Hf��s٘q��܃$Y�ဪ�`?b���1���`H���:E��[�&Ĉ��I��I�pt�c
`��Sw���Z>3��Gth�+����`��~,����7������TFw���/��ƞI$R�O������P��V/�������ސ��ޱM��'���mv@W�#`�A^���~Q�!��1��t���r�l��n0��<p����c�[��op��E3�98���a\:~[�7PG�*���D�Ԭ���sue���NDm ���TH����ș�1��:.�����<�fq����s,F�P���
��kO.�oGi�!����%R�s�[�c�~tK� �������g�v���[�uہ/X�T=����K>z����4�v<	�c��#�4�2?�:����x/�g��V�<O�#UK� ��v '���)4#�ږ3��Qf����Q���]f�䎡wH}�^*���2���(��s�
ն�`ڻ7E�	ڴP��蜼<�4����)�} �T��P�!C�	;r����cH�᳗�$'�|���s�BT\�'ˌ�ټK�����S�ȬC!���9�o��2�TKGS�Y�j�+�R/�6�o2�h���Ey+I���[��� u�],��YQ(ࢿ�`T����~0�
����7�	Ξ	2���)>)[h�ڄgS����<�)��HZV�2�Z������J��]|P�wK������	A|��?O�>�=i�=󮏤�=u>?0V�ciDx�؀]vS���<���1wuܣ�X�y�ۯ�k����������b��pw:�ζ�]>#�(�F���.��M7p�>� d�ڤa��W��B�'�.�)k�Gj�;e��h�m�!'7z �̈�*
vS��Я�E MQ�X���i��d���e$��p�J�Q�lpwt���h���iS,��4�i�%�r�v�d�>3�6mt�	\JN�k���k뻆�r��y5��P���3�?�]�����X���G�� �9���H.u�\���� ���~HT���?>W,8�[��vR�e2�|P��+(b1=lh���q�,�0q}h�Zv�Nh��݂�%A��2�yDq�A7cu 7ɮw���ϨLu�7���P���$�3��LI�
�?��Ų�TN�o�MN�U�O0�k�O�Gb��I�L�D���Qv�=��C�<KŹ*+��=E�2�h|��N��%$��rQTRE�����>>	ڵ�ۭ��O�]�82V!������ ��{g��w
 ����|o��_F^Eㄡm9ǯ�^�k=��� �!<������'�*�v��}��>e3��n�T`e���Կ�M�p��z�r�m@��8MV8[���������E��'D㊄����4��*{T�<�$a��e���r�z�p�RvHZQk��ޚ�@�L�������J��K�Y.	tji;Z��s��a/5���C6��z*X/aH��%�p���t��F�)F �b���mEP�F��~�ȑ�ʻZvH�j;�ݮ�Ã�U��Ê�O�*�ڢ2���+h\V��?|!�M�8}�=�)q^�@Z�8��H�IF�f�b������r~�c���[dU�|\�����s,��K� .Id.2��2���$S����D��7F% �&&�dy�*�u�)����l�*�U�2���?R��Ga��[v���z���*o�$z�F�dO+^pGZ���Jp�r�:M���sp��Ch��4v�r����b"$���[�s\����ֺ�����G��ɂ�6�)���=㹅 ��	��[�2�4���T�����0�㞦"6�S�3�*��g�������6���z"�ʍ���<|޿4�+IN�0����6)�WW��#�dΝ�5���D/MSez��vG�b��ėI��V�aЃ������/��0nb��|q@�Q{�ܻJ��}I(����Z��5 ���*?��[�f����bw�?-������͹���r7�Ԅtci�ى�p.��O�U��za��O���J���<�f��M�1|�t���ϱ3x4'(��,~g�<��~�H]E�$�aӿ���N[�sU*|c�u���n��}�!��k�kEC�8�S��������1Y�{U[��iK��뮬�r �	��W����3z?\v�稘�O���.J��!�bd�ϗ���,����	������B�&yO��K�D�>��>K)}7>�MO�Jd�B��i˚VG�ަy�1��ׁ��$X~�|���
�B>�)P7*]�>�����|lU��/)�Ty��}��R?���VCĹj,T�dOw��P�zK�`K����4ȁ7#�Oc�0V��8A��8�M�\5L\��,��0�=j2�ۨ�FO��,0b�`^v�pȫ�rg��
�)*�I��[�k���Ļ�������Yt2�@�ː�
$�q������Jy��N3���ػM���+k�u��,}��CuR٥c��I���-P����e�h�Յ��N�t8^|K���0N*1�fT��F75g���&�vCbg�/�e�����"h��P�)l�k���1Ew�c�n|�HZ�3jcw���Kb��嗔dRŨ	��2Oݣ�� ~��R��R�~����W�bz8��x���4T)0O7��I�3�,��*����_aK����j_�����7s�JTm2.Zؚm�ǎP�Q~�52p|U�3�9_��и>;�6�$�}sT�f����b;7�J;���Ώēn�s �.f3��
$�kۋ� ������?)��&���q`.R���"oᙻ����ٿ~�)��������?���'������$ߑ�>�f�p�}[�0+�7�@�����M�G�e�q�%���n�C/?U��Z�W��5L��}>~�P�=J���yBw۱�g�EL�]�,�0���}�J���qo�Qr��踑�����S>x8� �2|Սm*����U�MT��Bߥ6���z�!U�������J$>�{H�,�K�%g�{r���`���f7�,�"� ��A�&Ŝ���ԯkKbF_øڕ�ߐ$C��,�1��&�;�mx#j��Y.�c�N�䞄CF�n�{���ĕ:�(�ū����]�Q'��\�]�Ƞ�9�ױ��P{��Ǎ��C��\�ŵ��^ת������¦�hciu�(O�Aã�W[M�E`h�#x�F
�������4_�&��ʦM���(����S|�
���x�����i���Y�t o\���>U6^���. c��}�6���7 S�4_�K��S�G2��b����ε�TKp�XZ���t��/��n�6��6b4�f��)�z�:�j��~��1��<Q�����v�6ΪL�d*�����S����R^`��l�|+�`S�ܹ\5P���fIAJ����P��=0b��=�Z+�R��Kf�q�������r�h4���R�l��~�E��)�Z�@Jd�x(de��ޠ�ƨ��:�!��,�;�` �����>��Ѵ"U�\�g��@��]P���\<to�{Z�Z��L�<x�aY� �$i~
��+I��{���b;��,QAvR��w��	�r!'���E]PE�]���}	�?!T,�"Z{��uX��ٰW�;
b��x�it���� x��)3���+lVoiw��.Ymbu�����D
�i��=��0N-Z�s>���=Lg 'N�LP�2�ڻ�	�;��G�D�hR�O�kd�d�%�{��ⷺ�󝩁E�X?��F�P-���XKAQ?�KU��A'�O�wB�@�6�qK�1
�9��CG�*}���k�����4�����y^�8?ŝ!�4u��P�|{�L�遾�TU��%Q�Ԣe1�/�B6��R��U�A�*���3���OZ��]�u�9������ђ���H�.|Ҏ`F4۔!�zˁ3OOrZv�]?y�S~��I�
������O�ϫӔQG8��Q�l���I�H������v�[W.IB�<ͤ��u��>��y�8
%�p����f���?��^��E��� d{�3|P�Ǌ�4P�G����8i|������L�a|����)K1ñ�U]�V��_�_*-W�y�K��&|0��9�@���۴O��x(#��n!{��շW����pG�z[sJs~O�1j�r-/�o����vr�w"��`w7�����f2���w�����ք�/�:
S��kB�J��>:>Eh�T2_E6���?op��?5GYx�&��6P^���]����_`�4�v�q��+a����Im �.H��t㶕2U����5g>!�` �
������i��ޕ����Y��_wTM�Җ����B���G|0���f�X�A@�>�I�<���]�bu�-���X'��<7R���4/AG������#���Z���]�"�`�n���[�S�b�@q��,��'�z:X�`N<o ��F����`��o��c,�=�悐]��)'�:C�rB��w�WA$R���!f��S�Zpy�vUr�Rޱ�j��Ik����Q`I�(j,��-�.��g��D��� �L[!.�3�k�;p}��5S�Χ�CZ{�x ��R\�b]������v�u��܏�[ì:��P����bq�V�C�L�6o��q�u��%:q\(�'��:��%�h�j2��F��Ӵ���+�iOk�:p�Ct-��7]L��`R�YSŊ	{ÆlM�y$�j1����|_|9�� ��n�!oIeT�/�aT
���H�*�\ܠfi/¾��q�\� 41�s��1�pa~H�$�<Se�=x1�h���E�;G�A���j��S���Ӱ�~i,y�[���p��:]�1*��F8��A�b|�`��f#��mN5N�+Ҍѧ��l�V���)��Bǿg�B���h����iu*��J�kѪg>�o�FJJ��sh�'����,}����p�����!�3��^�G�ц��si�}X���1��є���»����_�Ϫ�1��ΥT�?�1	�*�f�'�P�Zi\JIm�[� �%jz���6��2~ մ&���S=��|�"ym�j��_3+��|1t- ��h/��@�#�����p/���2p�
�;����=
�Z��I��.@I����&?�m�	��"P��;e��ʨ�LDq	�$!b�������Snz}�Z��9���R�v��c�.ؔt`��"#:i����6C��ou�iJ��Ddxm�A�"��	��YY~0)ۧxϫ#� �m�������Ӌ%m��,y�$�ħN�K�vd�Ѡ�I����	TD�;ux�T�{�|kUޫ\*���+IaXg �Lc%�ƭ��� ������%#[i"����_�#�8* �!@Lg5� �D��*a�q6>M�a~���U
䀣���7��J��B��g��5n��H��~Y>P�W�)��Ce��c:1u8���ׄ�s��:��yL�XE��A
b���'z]姥�8B�����d܎�#�B2��ơ
U�3���4LT�|���ˆ��Y� N��賈
*�p�x�r�!��²�,Q�[��5g������?}�b3[֍P�z������GFC�#�[�������ZQ5��X���Dsy��qObjM;p��&�'�����A�*�~� ]�Yi�&�_�����
����j�:���2��(��1���c�ȬO�@1dR҃%��nU�qe�.��|�`J����ã�N��v�R��[q6�,�p�%m�d�mF�$?���$�?ׄ]ј���Py�����n� .��1P'�
�B(���4/�N!����l� v� =O�0�ul4�Q׼-=6a[A�8��"M�;F��!tch\z<����W�zs���K�N.�A:�i6 �	(r�k�v6�J�Y&��I�:��%?���$���W���d�J����$���Ak��!��͚=����(m��mT��Pþ�{�Câ-b�M�M��9n�E��r��x56/#`'rEbof�H�Z��F!����ǻ�D����ES�3���{��9e[;�W�͉�lL곁���e�'���P��֏<�Rg����K�	/:��.�#��AW׏����D��-�C]Д1 i��.4ȟ�?�a�!و�r�s���*�_����ٰ�5��a7��(����X�������=�sy���*��c�����,�)���8C��Қ}�>���|��mg����8����2t��ԧ����M���.�G�����b�b�?�M3� ֿ���
F��r�|�N�Η�m�Բ��l��Ѯ=c� ȭ:s���b��:
��j�n�u��u5f0�PP�9B���hh|�`�Rq��u ޟ"bz_�p�b��֭�4	h͋uG��U�d��a"[B�E�.�R��N�͵a�|�=���- �j�3\�������9(DZ�)��3�#�G�><.�����	l�6��N��%`�qٴ	j�v��]�n�@+Ab)���&vB�����iߛ&�4ݽxh�^�k���i���|�Z�޹a�ͅ���G��2������&@��K�(�u@%�r��L�T4@4�fH�T�b$�x��R�e�E(h5���7�Ԏ�"C��'r!ZM8�] �Z���,�����,HT�lJ������"���uqm��>ɒ�����f��=dKΧp5c箚Q��G$��s��e]ҩ��Ą�H:�d���78�H�-�u\̇Z55�w�*A�H*�j�
i���o_��TodVL�0_�r�*.=�z�Y@����g�t?C���0�(�6�V���8��'�Eܲt����˫-���ڸXb>cC���d�����y��)¢q ��8�و�i�,��é�~�n�}�3\X�=��:j܂�ԣ/y�b7�dɔ��1�i�z��<T�N��v]j�1¢̷XG��#a��@�r��!,G��5����e�:�#���_��5��<C`��fd{Bo�aƓg��K�"� ���bl���+��!�*��ʤ�%�k<�����ǥ�S�L���A�������B���H!&\q�5A��D�k�w�nt9R�[x%S����0�̑퐆�ƔNÚ��
c�U����4m#b����[R���.A�r�0�9&�"��]VS|�3�[�NIu��S�R�صcs�^8o[����4FsD(>�D�XtrA��p�����'�H�P$Is�`�>��� ��3���¾���n�d@\N�{��s�<�� g�����5��E��ŏ:]�С�ڑ�����1�l����@0�j���\m�y"����˦
 �"39km�!!��5Nm"�Gym������>9��]l�Z�ڴ�Ɩ�~C��p��1�?�B�VO5�&]�I�#�p�ZUÊ�} �iTj��,jX�~���D��� )��#U�Q�oڏ"g��`:���T��uo�~�qͦm$�0{q"uE���Ad'�FCߢ�6U|#9���)�ǻ��b�[������@����`sO�>���A4Z���gB��Ѓ����g�c���B�b��:W��hU���������P�����q#:2�3Y����3Z�(}c�I��W,B<�����N,�����־V����Q���}y�V�n��X;�N�Ŀӈ�Λ�żW��ǘ�Ȇ�t����P O.�F&+{+GH�n��e��	D�Rr����-�{U��x���� ��
�Y�4�Հ��|%���Y����eh�^X����Y�M�0���'�����"��Х����8J�"�)/��-eaɈf���@@�dnH�s�H/2�x��eq��C�p-\�#���4������PoqH�Aaoۊ�*��H��{�M�����1�<5�c@1��5O~��װf^��Q[�F��[Q�F1�%9}'���[��W����'���5	HuK���Q/ 8��T:;�{�(C��)��j0����)F���j󌤥.#}�&[>s�Q���Ζ�������6{� �s~�p	��o(ia�(-l��%���w�DF	3v�Ʊ-�0��]W�<j��R?�����r���N�]����͹7����1 �4���w���-��!?���?5�Ŵu��_�m���\&ˮ�>��q_?7#��<�j@�;���?-���򠆌��I�E(N��e��qx��QӇ2Q�&�Ϳ,�iZ�2R�P���!t1&���[��l�i�3���mA�����$����b,,th0�����'�k����]fm��*���!���籕SĉKJ3��Y]h���aq>򥉪�A�d`�	�d �����������86�d.CAf�
m~l�7��O*�wvbDap�#hH~R�4`2�Z�+�K}�L,��j����	��q��H�&��y8lj��-����� ^���>�m��1Amձ$�_�f�����H��ލqΑ�~�N��G��eɰrf���^�����!���~&�̛8`���! p�a�
�}� �͌���eLQ��y����(Y�p��	ncv�oa
&�.�(��J�2"�gѪ<�?<��-��z��"�r�!Fe����a��/��)�"^�ە>�R�9"ver5r|
�(!���K�[ꤖ���� ̓�������˿٩�s]�.VZ5��7����������&j�ˉ��.c2�X��d*���kc�M��6����zpe�F�x� t�j���6u��y��,V�Ą�a���K�h��Vic�//�t��E����S�x������%��<k�rJ�V��[�N/���,�Xĭ~���PC��De��efu�%���M4����o��Z�wq>*<G��f�_lђۣ�:�
Y���tF���+3�d<��*�IP�`����^�ۡw����`>$��x���D�+�d�4��h�7�F=;�8����띊E�	�Ī�m�oh���,���΄:^�z�&�Zԏw��;�
�pW�������u�<a�$e�T�O�j������H�;(H�l�����A��ֺ~5�,���A�5E�3���1(�s��m� �7�Y~Α�3h�pe8 -��Hh�uH���B�[x�Z����H�v���roT��xV�A�{.0�����e��g�0��ʈ�/����w ����8��nو�p��|ł=�I��b�[p�ε�?�L��~p2����L�u�ʼa~��$q{�G�cހ�g��AMl�}��j�bo�]䋢(�p�G�F�s��h����DA���]6���f$C��,�n��CW�7��N0^+��!������5� ��/�C�[r+_k0�:x���2��P6��	S�>7p��6��9�ROֶ�h;m]�/�9���+�&��BĂ'wӒ��>e�)O��*�l��c5�[��[�Mo��C�q m���|��g������̈�����P|"�)E����zmw��6�V���x������M�p$=�w��9��*�.y-�f|.�M*�tNkIp�7�#Q��%P��~�d�����SA�A��!���D��T/Vf;_�qyH<�|�eA��zR�J����� |�u��!8Tf���BqmL��3/���1̓���@ʱ$s<q\(�.�{����b��6[��F�E�院�����M�?f��42�t�\]�k
�k���z�LE[섩��j0؁����"�����U��f�w��ܱw	��tlD@�]��Y��eOg�ܭ9.0n1LnA�;>D�U+���A�s� `bI�ٽ����Kj���sx]�V\r��Z��-�x�����]P7�5ŏ��Ʒ������ߌ�]�Spެi��H�{6��+����I��~�K4���M���M�����Mm��ӆ�opK�G��I��d�r�:�`���>�	N��5���6;.��>#4-9�	��`��9���?�8�	y�1I,�%!�4}_DE��wI�e��5ŰO�OI�߁ iK=;o��c�sl����\4$%*��B�0���K�eOi�!bk �k���z����I�t�\�$�ȼ�\#� @b;�u��u��R3mW����*y:[R6��4dIb;�'$�����ȿ���!��*��1��wM�'��
�)/9� �u4$���g�Xz�s�>2u��H#W�����]�)���g2o=����;�����&�i����	��l�ڻ�HY~r1&�p�g����!z�̎{i<��A��*+n�N�7f^��{�#�sCQ��W����	Vfc��.���f��-+��Ǯ��{�i"	�-�Dw��X��x� �B}�xU��u�(z֜�Ț\����%���?��|�H+���F�p���c��c��M͋I)w�;{��TE�Y��`��;t���E��`�{����>�}�vR��8`�/wv��tO"���|U��a��BH��/>4m�2�2!�t�t��p����Lٛ�o�]Vk:8�\4S��)Z�3��[��BL	Bpк>>��S���}D�]�y!��E?�PR��[��//���t5�b��7@4%��K��b� R�]��^�`m��j���<�Ai9x���w\N�F)n���({�,L+l  E&����Ԥ�Yv9�F]oT
�3�d�f��W�xN�v�>h)N6��h�����Qz�/�5(&OT~Et�t8�D�wK�=DA��e�"�?a$3c��փ���[J+ ��6.�j�R).P�u�Z>,��50\@)��ݲ�5�����:�R�v���9�<�Kq;k�z	^�oo�Z"�`&WM��c�sｺ��0���uX��-OɁD�T�R*T�ޠ!Ɖ]|ӬR�㟠N�78�!�����*2K��`��$n4�2	�b�It���W�<���F^W[њ,�2����B@��;�R�J�����,I7\�ܺ�i�w_�n|'��*
�!���Fq�}D�09�@R����Dڠ&�� ���	앿��d'���/�L�]���b�n�\-�٤���$(ϥ�A�X7$�n�5� �lk���YP����{u�E��al��áJwi3��dB�e�b$���9D%����8�&���7���:����Q�'D�U��k7.<���D���hz���J/���?[n<�I.�����<4�����}�q���s�Q
|��D�X|a1�E�sIn�h����^6ۣ��M��Q���%�Z���4O�NH��kL�y)A�	|�l�lA�E��i��˝�2����q+7��᜽,ejx�՟Hk�󗀫\y�C��;�ܓ�1j���nP��Z��ݒ�������]��bb�A��5,15�X�it������$k�Q�o�Z��Ix.��&I��u3?j��q+g�Mzz��X�z�mAe�Q����[a&�Ǹn���u`[و�JV[��t3��*�]<��X�c��������اJ�i����E����)��n+�VX~��sb[@�R����)c���y�#�����gD���p���b�5�_r�⩘���E���"(�O&E��3��K�N�c(&3^ k4�,rm��Q���oCe[�� ���o�;�-�t�E��+�,��"yմN�,��~g߱$�=�u�������!��|�'��V$��J�4�(���I���P}�b+��(jr0������W�J�eCQH��l|����Mm4�43�rY0J�:D ��
C�{a�%dls�Hܯ-|�l �b�a��}+�\��ǥ�<�Y����7��&b���3�PB��}3M������,Z����f�k��6�����@��ߕmy�QD���V")Q/��w�+EP[>�jB�N;���4j�Z�YFKYi���N�jNB���	�C�-������^�0T�1_y�K{4��=�ݙ�ӱD�WxF���lHd���y(�݇�2(َ�梎NP�O�? 8��w��P��Hu�eDު�����{��~ ! ����u0̤cR`%�',Ur&dZ{����	*$�WJI��a\���}mړjl�>�){��A�ik�%��D^��P�i�Lr�VyX22!&����8�T�.�`_�\F�8��_��p���a��,���(�؞������8I��[_�e�E��l#���d]�7Je���_/t���:q��ȧ�U�o�W��JJ�p"���fh�B�tx����e�:4�#��/b��:W5L�O <u�Ϗ#;#�h�+����	I3/�9�Kj����y��4���:�c�8�n��(}9��v��~34W�_W}�6�Wz(S�������M?��L�HDP�xA	>
]���j��%X��퓒�=�P�L��Y�6K&y��F�;D���zDtI�`�,\�Eu��:�h��aBZMN��1�*�	U~������pp�T�_k�9!��V�:>���N\Z#��{ ���W$�i�ϋ�����ZK��P�%6�w2A��x~�1�$'2��L�/5�b�U�O>�ce~+�H��)�oF��(r��'T�0��]��V���,_|dK�.M}��&�!C.W�Z*h/�qi����_2+d�Hy�����0u�K�$����N��%�Ǣ���eT~�����3�*�b�/���蘀��W&g(� 6V��SŴ[�ק���䃵����v,ޢ�Lz���!�H2���g\n1!�D��7z*OӻЍfM��~�K�m��Џ���So��P��=���l��O�C�� ��q?,����FPj���@�%[�M�v߮�� X#��9q��WW��_�qYF4�jk��#�̹ɽC� r[h�㬰3�J�.;Š�c�uW:��ޡ+(�l7� ,��c�(�~e���W��桋��Y6rr�6B���!q~6v`��y����.is��0*S��-�0�U�V(����P�\����gay����1� +��z���d��)������gx��뢚��'a���F$�����+�o���Ԁ0u$�.6ǎ�,��a'��{;�#WA���RU7*p�k,��h�[��u�S������zvL�5� �rg�5?ґ�8{N����w��W�>tگ|�P��g x��G����Q2���$z�f���@Z>����@��j������[7��qI�سq�b��5�g�>����#�P���r)
>\���Kw�Ջ��|�h���Zۋ���7q#�:�s
9��5�j��4�g�(��h�����>~����ӯ����:�s��Ќ�豀�r��=|ֵyS6�-R31�81�t|}Z�C�]68l�Fs�<��AV�L�0b��>a��g2&n���nf��B�"�h�q�6�k����iJ��Bi�]R�@� 	��k��BL��^�ۭ�o���:���KfQ��s�n������ ����v��~��;�������D"��bQ_�{�R�^�Jϴ�|�젊�6^�y`��i 	+p�0"ZH�fMSӚ�	K:���"�Y>Ys�Qq��]�S��)]������r����GA�W�������0�Pg����� ԴG�1wCN8�1�����gO~9�]���{9�8W
���w٠__�N��K��E��f�;�
�Y�܏K�aTjoY��!e�D�<����T�g�!eg�IVn*���d���oxF�̭�OwZ1!Ӈ��hPhW�mł��4H^ng"r1��_׽�(W^tL~��W9iJ�b��c����$���{v���f�.jzC\��\��nW �� ��|�щ	;�I���|�/���=Ɯ|�62NM�i�� {�6Ν�wEwC����߾�Nłz�v�en�ȕ)�8��F�3��Ƒ7��BX���'�H��Dܘ����:Eײ�!�LX��j^F���	MB��ꆨ�g��{�������Ȃ�y�#�_�'��Ij��u��p��z����͙�%��U1��q�"�hue��A3�1x5��q*��Z�����g
�F����ʖ��!�~��^=��ZU�L�������2RX5p��$�a[>�ĐG6��VCKFt>|�<c.�L��/[�<�e��h�W��utI8����TG"�����
�Y9vӴΖuf��$��g$��!�V��G��4(g砝rr�?2�e�Ϟ��x'`A�����������v�q7|�^\�<��-������\H�!����R��yG�������(�vSh��e9k1n6�� H��k:*���u�`���>��]/�lf7�r65����3'N�>���@#�9{��|Kd1�T�n)��U񢐽YL7�:�p�G�j{xp�<�ד�t��#�Ws���Z��A��5���{��bo��H�ΰK����N��vQ�<#s��3l�>��GӨ�D����t����P��*��c�JՑ{����Y3���{���:�㝔�7`�-��q=ۚ3xF|����|U%����\�[�(Q��6!��m�x��9�[�m�2 #}@Z[�"B�)iK���%ѡ>{�3�q���S�a^�I��+h+�*3f�#��F�T��_��H��jpm��`O�ʒ�zY�߾��Nv���(��F���R:�q8��>6�Ģa��q�����>�Q��\ro,i>Q��^-5@N�����
�>8��J]�"�|cŊ��==떬���Fՙ�S1)yM��F��[�0o�t[wG���qv�4��|�@8i��.lU�a�;|�����1#�]��t16�sOG�Ќ��t����vj��Weϰ�H��ǽ�DVve����J��6���ߗ?Lˌ���\��M:���S#�s 6!H�֏|��S,��P)'Fwd�}	��99��<��ڃ��4�v3�!���^8웝��m5N"��n<,����_1�-��;����mѭ/�l�^N��r��hJVsᒳ#qe	�ԑ�����Ψ�Ns�5ֻ&W�F��狗V�D?㫼���/�*��("�x;����X�t� �g|��D���b��>�DfT�&���|�����o�/�P�k��[Ԛxd�H|��W���W[��n���t��x�x�e������c�)��rh�ÿ	��|}26�EG���g-a6Z�Gkj&G1	�������t��2OM�h����w2*��v�5y�SK�{�N�\��!b�L��I�Ő.�&��
M|n��eնmt�uL��>w	�ɸK��G�c�k�DҕLr�A���Xke���=D���%�[m0�_E�0�]�x?~`���V̷MQ�"O0a�i��,���GA�.s@�ha	o����|���-��&�{el�؎!��|E�U�Y�^F�>���q����	\����
ÀC�6���]�+���=�lq���Ύ���\@�#tU�,�� z��DKԿ��yD(�.����*o�ǵ/:!M�<�6�Y�k�/3���'�-&�&��z���KϐNV9E{�_ �lz>�Ka�<Ra��B�h���!��v�w��A��7��)˨Ĕh�������E�Ͼ(7��mP�"4b�`�<A�/:�TE�g7�*��`'�%��u*ƿ~#xr^�N���}�"�b�h�$^d_�l-�-�]�!x�i'���3�hjci͓p�K�9�ұHqr��I3v^�}{*�<�"�W�XnM�m;���f��(�H�૞@�{�;��l��� vS<��N˺rq�� _j>�ܼ�oPsĨ�=6d$���VޙhAs�b܎=� ����u��pA�1�d�b3�˼:��xBƖ�����$����ʰ]����Vho
־��Y=��5�Zݸ���}QƋ��]��һo�"��,~ ���Q1�2mn�D%/o1���*g�K!��b�&���A��B��I���Q�k�#9�;��p���=�پH�@\�����/7T�?N��sp���k���w������_BT��sW�܇�%ʦ%��ԹF]Uqa�f��~'*O�k�|L�f5��*��k��QjE��:���^�����[������S72����r�p�T�k��Șu�Ow\=�X��4joq�'i�g]�)�X����0��Ʒ�\5�5�9�o��>wLy�6.fd"���~�O+��`<"�����Y#UڬS 4ItaE��K�9M*�1zu�Ѕ���&�G݆��öe�=��z���{�8�f�;��%�	$�x;|.�,Q�
���TQ�mq�$~��ъ��}�ϕ`4�^��5h.�H����v-p`��eagNo#X�xE���)��ן�7�U��8-�芁���K��^s���R�!�O�.�n��N�B���`M��$��h����[�?�_��?,A�3�\E��|@,�X��m@��X�m��t;@E�̶ -��R��U߮�q(�(�O��k��l�ZkB��a'�*b�9��a�����1�3�+ջDc��W�0��:�����5)LZ��1�R�i<��\�U��X��7��ܒ{c�܎��E������y.J�Z5?�Q�T�Qŗ�,�@VXϦ`�Rmk��f`�`~N���CkϚ���Oħ��Mmg��vGc�����JnF���t�.�x��y��mp�W��Y��̵|���zj�\�������sf�/XX$���^5L슲r!oS�SM��ˀ��Hů��>y�cA㍴Ԁ��k��0he�骪��3)����؎��ݶ�-��$��߼�l��LV,���z��O�`��2��B'�J=O��������^"�i�E�)���Ԙ��^��f�b;KzWxo7
7\b�$�dmϤ0L4?[בw@�e�ڱ7�J*�%���sɝ/�Ŀ�Âй��*�N�.�5*xVXƙ�Xpd�&��gA�bnc�ZK��Z�!@e�!�{10�vA`5���`�9�Ҡ�v��H�(�0�8���ᕴ�eBJ��Ci�6$���.%[q;
$�w�0 �"������$�����C�ƽk�U��\H3qg%'��K?ۏ6f'u�M�T�M�7i�C͢�>c;���3�ޘ �,Ή�&�A./����`JGx5��հr���)��[r��ř��̲�C.m���|��V�q�ϬܸK]9=���b5�x,�:Q[�K(��j'�Z�/ �4)���$J�!5yn����o�D��m{oЍV����n�xJn֕#;��S�#G���tq +��՟�^�{�n��Rf��ڛM����r���;��q�Kj G��k���_ϯFd���0�k�;9rmH����;R��♮�!``���\����PGiI X�(�T1��<�.X�TR�'�̌�>P��8$~��Y��%}���0xS��9���j��@��w�LȐ��P���Y:�[���s��vol��D�H�:K�k�:l��v\��s��~+D��2�����3~yّ<��.���P�A}�o�!b��RݻP�\���Wf��a4BۇFy��O_c�nH򇂐�A�o#�� V�&�-����=��L��y�:���,Z�L�̛�JeA1�I-�K��׹9�˪�+����  ��1ٵo��w�e��ǥ��c�d��j��pdII�>�Y��5����P!��e멺iҁ���]�a��Ź#��H�4�_�0�X�(�jI�oz�U`R�`�D�|w�\B�q�'����G�'��\��s�P�7zɔO��򡈥`2�5�X�Uk�����B\�_����+8, �f��&}G����t��ٚ�����d-	��a��ʨt˰�7���gW\�l�_�>�!�f\��륥܀����8A�2�χ�R6C�Isy�MX�5j�x��2̲��t"�o��nLv/]ZԼ 3Q�{��#�H��ot�i�%J��-����q3+ϓ���P<��.��"%�U�r]�)]��>�}��i�=q�"9��>@���Swƨs�i�%T!�C�`f]�ƕJ����쀌�������g +�/�ρ�f�?��j�ؗb>h��k�`��.*7�*��o�
P��|�?��B���b�޶�Px�浛�u�%�%O���&��(�J�L��`!{��r7(تJ+[k���Sfn-x[暠�fab����:��$��o4l��йpX����-#�Q�JJ��6ۢE1�C��c�"�M榧_+L�p�����`@C���^?���)�{ �:��y����%,F�O4(�eZנ�����_6I�H��q@�Uso�\���k)x�z��Q�$nfS1�r�V�0����2�1�SqyX�ƛ��p<�􏄎k���`�Vg��=�ػ~�vy�g�
!STT�K�]}�I;nm�>w��1�TQ�3k�r�,\�qq�엌�D��&.��;̹���9��uX�c��ЫLP��W����U�ƴ�'#�OL�I�3y�I!���)��k�w�$ά��D�BXNl�(;�T�.�j�m!�m��-���$T��~�k;da���-��8���Z�2ͺ�2}��1��D$�I9�"�3( C��S�1
��lt%�E��[�T(�sݵ\�A�Y�[M��Ia"p3xޝ"RYch�y�ټ��V��=����r�E��%D00l���:W��0��+"x�#���,�zpK��Z�^Ș������(��$[�x���G!Q����kg:z���PR�����F��������L�GQЩ0��r9�&)�0t�����/��d� ��M
]@�Ѕe�|!�;)����|H%ME��8�YF	޴L�u- r9���t|hy��KZ�B%Yķ���T~�ޣbKpJ�"�_��U�}�2���"����}���W�va���~J8S�$^���HXˡs�U�W����at8�A���\zU�W�'Is$"5�G:nu��g�NOw����B���?�����蒉��d��`_в��)<�k�kQ�q��� ��u�j%Z�@Ļa�u�A|�%�eGSnŸp2�{�'�'��<e������0�Z1�L�xg�m�&T&<��}����qX7�%% �Fy�[�~���]!W��&���
c#^�/y0M��ʫ����>tB�F:��3~�'�`/ɜڿ4�<0�j�ڹ.E�SGX^���+5k�p���h}���ث���0u�Iv4���#����tJ3I��L��+�c�>�>�9�g�龜�����'��號�}<^x ��y��z��R���q\�cS�d�2�U
�0�2FJ5O:N
���<>y�l��_?!�T��|�lR�')����4�x��ju��jR%;�XӶm��$4��T�g�+y;[�l���P+Y�~kg��K� N�`���V���3�B�����^v���*��*֏.�!�ד#����b�
�1����L�/��'�RW��S�:a��O�5��f���$A�w���U� ����m��vƿ+����4oP�f�F*Z>�����J�O c﮲."����کCy̤w8�9qT[����fCG�`N>�x�<�C�>�����5�;���u`C�?<�-3����h�@�*Ԅ��6*���-|ww���{�.%hT�U������Z�,�����_E�@����5Y��3��֯'mMs9�@�]8⍍�P�f��5M'����d}U�P�E�(1
2>�"B��`��O�ly�t��q��Gɦ�OJ�*?���*��B[�53�粌n�F�䘴̓5u��C�m�+gis�e�|r᭣%c��d�r㣸�#Eh��E2Q�\cN	D��� �4cf���Mշ�3��k��6��y��!���D-GE0;��0�&�������O�L5*f܏n�7�=1H�f�{%ܘ��R�y��Y�ӔO�����\2~h+���x��[�q�����M�^�φҳg9{t3�0Z��~;y�p?�	���@��6#��i�z3�K?u����>~~qm�������k_��WH�c.l�yA3<7xS��2�Uό�]8�f;G�r� 2W+햨��B]i
V�i� 0;�ӌ7��{����DѧE��:נӳ���&�����<��Q�ܫ��cc�1��N���Aʔ@�U��Z�A��V���gp,Z��F:CZy��;-4t���FքK�Zi�-�1}Wm�{S��d����{��+tXfr��m0]� Q#�x���V�����W�w$�`���K@���$�H��Nn͑I�M�G%��f/���7�JȯQ��G��\��J��/Pַ��+8�qR���<1t,���d5��U�m� $2�5����q��]T�{��/��R�GDl�,���n�ߚ��0S	����ޮ��.���O1"�l����[=2*�0�ػ�|��)��D�#4Xq7�^:�3O��D������~���ʹ�~j��v���0�E���=��D��$��j{��5�o&�NEYf�Asc��V����߇Qc�t��b@�R���j�G���p�`�O6b��.��OY�1ڤ�>��I�`������Z����Z�a t��Cf�l\�
�pe���$�{��y�O��v�|{$#��d���������^?g]ˀ(���ʗ��"O�?U�H���+�T��IN7`a��p~��.E�LM!j��Dث��
9�#&qZ>���|~���Mآ	�H�d�W�*�SM���HL��8(�Jo;�����A��P��;��tt��c�N��4��M����fP>
��K�H�.�[�
D� *Ţ���{Hc�(� �~-c����_�L�����J�o�|!��~q�_���=�'��w/��k�|x�7�\���<=�J�~�]�f�LVGL�;��i_.�G�MԼ���#�ǣ��Z_XF�\
U�U�<�p��kղ�G��)�SJ���P���z�: +�Z��r��9��m�4Z�:{��H�_�$"��<�{�+��l̱R�E��9��c��D���(c�C'�b&�1l�2t�=���{�D�1 Z��d*��'E����N̴�1#��h�Ya���s�e���חE��o����jM�MRk������h�|w]m$�vBP��a��G���"=䏜�z���R\����b�_J��0R�o�$c#�
4�� �^�d�KDH�Yz�IH�(a]|=�������ᔇmmmG����䘈�H�A1ϙ��D�-��z�(�o՘��@�=u��dr��2���sCA�Ќ+	�9z��ik�1��Z��aΑ�V�^����.{�A��+��'�Fas��O��X�3O���)���T��A��w՘�5>�Ip{d3�V��� ��	�B�ep_aN����2 �J��:°��~Q�_&v�6��8[�V�H�G�e0)���\��z�w���d�W4�c墹-�/B��!�;��3��ei�N{ �`�Umj����.X6`�Cz�T�@��F�N9��(?��Eg
(O3<JM�~r���b��t��An���3��S��`O�t{�쑾�5E������Ԝ<e �=4�&�h�7������?E�;��p�f�����IU�؎3ٿ���-��-�`�ǀ�:^�2�\+��Ć��sB�G��#v�A�Q�"a�h��M�	�/�!��6�N��g��.��-��X�[o�ߗ��8�e),��l�>#`qp�kl\4���lH���U��N���̘�������P�!�b�J0F;
!c�.���S��G�U���X��=�7b��`�ua��9k婛�����,���jU��D���	>�kvU�oT�jS�i<[�p�q����i��Qz��qt�����D�/rJd�_\�j��a��N*0�?�|9��������j�J1��s�u�c�����P,=�8`����(�߰?��5����ވ�i�ʵ�ҷjc�����1 �]~�>�x�L�ERq7eO�֓@�<ԩ��ԚE]RO�߈��x�r�d?�J�͚�kl�7����Ł�����]&�uxy�>��9�w/]dN�f?���Tvp�d '���K�$ _�Z�FY
�6s�Ll��Ng��/�x��8����b�C��fY�p�Ԑ[��g���(k&�;�.�������ƈ$�IK���4�0Ye�
�=��#V�������(
Ѣ��7�;�Z=_�R��� ��h��[�*����.���&����d��D,�h#���!�-����1�ͮ�o#L����5���G��غ��H��r�k���ĵAm����+���r��A��	L�{�v�ف#�CT���,�Rƿ����~J�t@��/�a�ǉ������˹2�*�t�Ec:$�Rl�M�GP��%��kv���Yr}�~Y�ʾ��a�<�N8�~��ɭ,٬7N��J�UL���a��&�tChx2��B���켵�헬9�?�;��E��x]�y�bV��R�N9Oqa��]!J��S�#� g��C�p�?;�n�ѿ�8�sI5�Pǰ�/��C���]c��ӯ�4�eqkp�1���T��E%h�oFcN�N��ڱ����0h�1��]�I$��o�����B����0���7�e �>a�+m�D<��v���K�h��<"�;>��Fi���b���r�	H�5j��%h\IL�R1|�g%y����ͧ� 0�F�_�Wm��(k!��+���7 ]�h:�6];�8���Z�k��N+�s����DU��/�9�|_��֙���܋�}mYxAu8'�4pW�Ƥ�!Ft�th��1�����o��9�|@0��]��w��Z��/t�hK��'���o��:�T`k+"%ӭ�6�[���<�1g������Bu��sX̒��>�&�_O��xڇJ��+�:9����)e�!�S���#��C�ʘ��[�jF]F_��1���<2�ث}�d{�=3x�D�2��~�u$������=vh;�oR��-�6�&'%���oCѢ8���/4͖Al;kYz��*M`�HGF�S�V^�N��3�k*��b��3X�e��+B��b}�q����Q��\��@{?~��l?%��2û���3ܩ&ˡ&��Ȝđ�0x�{��T�T�IT���	s��<B�c5�<E�_=����[�ӑ���_oel�st���P�$xhUp��?د�'D�:m���;G?�ѥ2%�t5�/||���X:t,����l`��.���r�f8vyoj�v.eeJ�Fܕyh�g�N2`@Ӈ���5�d�Ԅ�A�S� n�^'2E��*�\�"	N�G�cux;O�ï�}�lА�2�Z��������D~��wPe��%N[��?xd�ʲ�`*�*�+�a��@�J���B=�\�Yn��)���}&�H���1���8� m
��2�i\��a
X�:�3[�����;	�m��"���7݆w3�Jf�7���CX)r_���X�@lɎ-� GK�}�$Fb2�b�=ҋ�`�]�*��I�B�}��Q��|��CP�=�G��B�Pp�u�k՝|,�|O}�C�G� wm�W�?xsn�n��p��L�u�kw���j2���c�-g�p"$�g�8�w�K��9�
�⁌ ў/�{�9��7r�,�o�H��s���:�Lڌ�Q�ve\�!��W��۰1i��y���nsbV��*R�%݊,'U���
hh�F�J��wϟ�9���F��^~<�^ �Fh*O�J���<���M��|;l��/�e0Ϗ���s�Y����
 ��)�Kn.��_1��z�`���[�ฃ��/��m��bW ��Yw���U;p���=s��W�k�+�jgkVb��Dٻ_�y�zFh���AX���%�G���;��!)��"l��Пf�2���
��,P�8KL�T�tEi���}�(��~��~b����v�o5�8�P�$f�d�7��#V�h!�����f���z��E�sJ@*���_a��
J`j�x��/GU��@���OG�z!����o@�9��G�wq�������"OB���o��P��e:��S/%�S�u%-k�M����WP#�?�v���v=�)��9�,w��pe�8���M]߿�a��,<T�u�?~0��?�*�p���\�>W�����L�l<:��
6,%��T�o���
߲��%9R����Z܉{J����<���6�_�q�[a�g��vW��b)ŊJ�')���ۂP�+���dc>3����	Tk�z�̘����1��ض�S���q��o�~��L�����<N���|�ް�	��3�"���<
A�]1��cDYj�y�`�9�F�K;��T9Ⴖv�]�)֐�zۍ�'�P�؁�z�i/�e�L&J���J��98K���5�i�{�w}!��'�z�b�b�3S̘�B��>;���	 ���N�T^�m_Ǡ�w
�8�$�ȟ+�-���Z6b`*�IA�@2�Q�ʿ�2�fb�yl���$��K��=��ZA�?����k��|�V �mt�m4���"���q���X)����eځe [w�s?b���v� Xſ��Ԋ����]�BՂ�)bu�l]]5�/0����"I��͵�2�8�L\u��߳]U6���x[�I��O㙒�Bg�/V���W�U�ub{�ơ���'���'ɯ!�J� 8Prā)"�����&�`��� �ĕU�M��h�Oz�!27��*�����*m�;̞N����Bu5to*Q��[�y�bn���
��y\Zփg�-m��n�:�PL##3-�nͲ�~��A��� nM1��s9��N��姏y+��E1ZZOm�"��4$��޵��A o[$.[��9z)�Bm=�2������N�Z� 'Ln��a��1d�����#|�X���}5{f@>1@KA;���9n�5��VEj`ؠw�^"ä��>D�5��;��� $}�F,>=�T 6������2�Ѻ��t���$z�j��͋��T�E/�Ó��57ok��Z�I:��u��D�D�3��(etX�a|H��a:G����%��yE
{��z cTO�.�{vƈ�~��	m�=�T�0*��C����1Khj�lk��,C���m?V�+0Y&����#�wwũ�дo�y��:A��7a�*���c2�ҩ�}�kO�]���H�H^r?t¥�et�r.p_�@��j��a�^����I<J����?3��A�ot�ǚ$�@c�?ڶ��O�}��ߐ��i���7�:\����ߵ
h�wˤ�\����7(��[C�0��cdW�Sm��{�[�����&r���އ�q*1�F訖���;��8�4���n�<s�n��H,�ᖯ��n�w�`��������Ղ��t��ȋ��!��;S�w�[%�c��|1�1�d�Ժ��$���{:�/��l)�����ޒ�iH�����������s��l�}�yc��Y�-޴��&��-�Jd���\~XZ��٬�O���,��=�ftT}�^]����ջ�"@?����j��_)�؞Hfss�|iT�="�1~	�vϮE�:C�;�Gn\MrzW-I��%]#��b� ���e"c>�kW�Ї��U_����䎂kT�����t�N$�����1��u�'��$�����ړc:�L����x�:�j�C�NKz������7 �m�Xؔ>�P���˃H�Ր�1�Rhs*	�#��M�4D	���g/k���dw.3}��;�d"�BAS��Z�Öt �sc�ŷ�7���Ce�����g�K+�=�_H��2V1,oc�'�#�
��)~)���lJ�?i�~s����s�ޔ�Q�Ř�\���[O��+I.-��8@�l,��!�s���	�?�iB��ޑ#�;�,
Y��ǂ9߃C�Zx,}�N�@�R(����t/N��*�Kq9���skw�Z4Hi����`���ؖ�!�w/YH�*�5ٵ4��)f��~�f��ebxաOgj�6�Y}���D�}�~?Si��(%+�U�����[���߻_�H1k��;������At܀x^|�	�Q&Q@�h��C)b��-�K�8,�n*�
>q}l�����J�L���;G(�s�R���@�V���2�Y�G��t��Na�r��$B]�F����;��A#��Ղ�BD������J kE�1�%b�ӶgL�f��¢U�kKY:�OѤ`s�K��r��iК���@s���*���´��wg-��:({�na/����w [������\d�*�#N�-P�ݛ���l��:!AY�l�F�NkӒ^q3 ���Wщ��r0����e�SX���mN�ҵ.�5�P�B�B�ȴxߧ͂>�?ث�4�lDq}r�$��h+_�R���/����Gg�()�f{P��.�i����X�sV��-��Ⱥ���vI�RJ��O.�C��p�%����1׫H�(;��ƀg�]OT>��X�b �	+G�*բ"0L�5����BT�~���"N�uCЅn��X�t��wc�T�fή,(T�7L����M��BMƞI�2{n�J2vB�o��۪Zo�ʒ�� �'��xL$�UtR�ꬆvzE���%(<+ʙ���k��F%����{6\t�1�s�N THed�2�=�E�i��.w��l?Y�%�ר�v���<��É�ky����VNRI�j�J�V�z`QN���_#'8��(�'�X���ˇ�BDm�uM$���m3H+���@P�u�s����~8��pv�,�e�;b"̉ƈ�'��m�0�ټP:����X��i�Z0��2�'��Ӯ]�J?�%5�m��T<�t���nw$�:�@�9����b�-�(�cx�)����>
}�DQ"W6czpn4~���)�sؒ�`����'�I����y";(���d��"�};#��2� �'BiH���vr�N�d�q}�$��Wr��1L-wm��̕��Z
��NQ��V8�5���v�ަǑ�od:��O���T0���ɱx�D��i��b�
R�g��Q�=[/�0��+�lF�2�Y��:'�P�?vg�����Ȏ]Ej:1����F��0SA�jN�N0�����V!�u(����~�p��fj��<5����G 
.����Bw����D}�3����]�\�6&�WX�/s�4�ȗH�-,l�lmP�'.���Bs!v�����9�S��/����j��S�7��$4��oǖ��)��U?�m�7�!!���:�;\�<T�Q�0Ag��a��%��ΰ������ZC�v�t�j�p��IIt��X]1�g���Mٵ���x���Pl��ql�e�nͻ��t�]��.y���
��(��	�~���NTr�h���V�y�6�/$�lAJ�Eԅ�@�Ұ�ȏq��;k�"�zi����_�����K?Zי.c"<�>���-�[U�^����=/�����ͷf�=Zy��L�{�R�OC�^�v+/Jq� !�s�ü���ys�@T'��/��S�Y�-ͅ�Y/m�o�.�g@������}D@�S[vP`5J��,WE�77o��K��J����ׄ����bT��r��cY�s��i�R��+�p�e����z�!.>_�A���=�)�o��rtWiz��.��Z�n��p�KB�/�f���:������[Wr��W!	G�\k��fv�@���
d3 ��D�h��v����~5j�+t(��zAr*!}Rxǻ/��罒,��E�R���������fo&8�f���^~4�"��Z}	h�mM��U��V��Zn=2��F��O���?�� V���v�S�|�f�u�Ĕ���_��PQI���>i>k7���7W)��
���ZSj�ď�^<⊌��݈�h��O����Uv!J5n�
~T[&�YQ���h�$�M�9�W �Fȿ�QJ[tr��ia��%KD}�S��&���wdt�&0�˴���ט�#�yg�Y�1P���%��Y�����127�8oqc�O�$�99���(����S=�0����^��9��fT�G[�V�]�cr?�E�=�_�1�R\#c��훎�qv�M�~S���	"���~3,�ϖ-�o�5��h��V�s�F%ZK���w#\�_�6��^�Fh��ň{V������.�rQ�fv�zw�������ݾ<
���$*��>�O�%�L'�F�f�n�UM�ׁS�0��,�!r�-J�%����+��.#"޸y�"�\�;T���skS��Qg�R�l���O�����gQ��2��$qb1����d���&S�|n#�\q�4(��f����r��	�3�W:�g*�gm!��U(�������^�u�F%��R��k�ҽƼ�bn����~���L�Kʣd"lP,���U�~�H��O��ȅߧ���}�)5�����8]�I��	��c�ե�8�"^z�o��j����`�Ko�gmF��tt�|`ӴZ��`8������n�Ҙk�����Ħ)Я��$(���n��"���kpѬ������/��exP���`�?�癮�̺*��B�A�oOs��H:|��vWe�2���f>��-��㗿��f`H� ��s
���K��\Y�f�t袻�ǚN�GB���eF�08�?��G@#��&�j�ϾM]У�#�P�+�=���8�޾����L�Fͤ�e��?��9Ȅ���
��~�&����)�<�+4���ꞗX�b���)Q^/�ڏtsa2{��؂F#\�D���uʦ��A��gMl�������4�����H���K\#J��\}�����&,ӌ����������4��z�6D��f�^rC���$��`��qe����h�Tu�ʑ'ݺ0"�(��?�L�-�\x���es��qA�Jwi�B��0M�F��xMF� �4��yr���{���N�L���y��U�L����W�r��$h�݆�UO!��gD
 K��t���C���S�}���Y�XU޹/?�0�Lq�6dK�LI<�&��Y�!�`�����w\],,'
����?�����뗶���$WF���'J��?s���~��@b�jc��`�#�}l~X�
JO���������@����E�z�=�"�t{�T�n4)�Yn[��{{���ع��1*�d2�{�����PD�gHa�:��tX��7j�v�&�K��ﰱ5D�öj�5��E}��~�E�������=���YO�`4h|,����.�}��ƻC��wտ=*��E͞���6�o��&�����h@�	 ����,��!������tP��FAj���FZrb�M������j�7���c$Y_��J�i�ųX�������#ώ5u�PP��Ԥ��Є ��	����c8?�"��i������dsv��a�a	J����V�Я�k�I5>M����h���Kp6��@�u2���@��
��%L�J� �ސG[ ���7J����a��y�hw�S[=L�6U�	I����&B7-�!=�R���L��S8BT@Q1�lڕ�"����R�>�zQ�R�>�]:�̻eP���/r\k�]L����yǅ��%u�^7�;7U������TsP�Qb����Qx䨼'�����H��B��M���H^@���ܢ�O�	\��ؔ -x]b���g^2u\S�Nz�(!�U��03NP4X*�ɴ��E�P�HҸ�j䁢�v3�û��xy�����[�zwu;��ٴD6)n`6H���h��n������Ժ�������G�04�	��1�M���f�|�t/-���<�e�����[#�!��Nդ���3q8���e�������R������,$8��w-�O͐�)mi��>u?�5t�IȾ�8.�K?�-1Q/�ux��d�`�A�m�$Z��#�5k_�?�|���ķ�8Q����}y��M���1w�
�
~a��5�v<X�ȵ�v���G������b�#դ4J��e��Q�a��Q
]l��� ��K�O��lCl*�- ���XLױ��ua�C��6����3��H�8g�ğ�!�v#V��w�?�&��o@C�U�g��m���Q�wuO���4�C<5�a<)��#�xl�y�I5�L�&��|m��a`�JNI������ư�8ս�s&{����|3y��t'��Z|��<�T���G9�mëT�-��ؒ��(�:FZq�Q���)5QT�
RA&�\��>�һe#�߿uZ��h7/��T�Aى��^��q��-w��J3UH���s4�PC^�3�[3�\�YsUL]�;�'������Y�N���[�S��U��0��h� Z�Re�����b�5w��A��� ^p_�ۋ�SfD �z̓b�S�焎�h�ߌ9�z!��@M�m�c�C�{��hzϤ4իW°M������	�E������"��s�။�$I�A��'g �#�R�����SR2�|f���d�N���q��*'P�/�#A,nQ(.<� �L����.���3��	��jS5��F�����Z��>VQ:aeJ����T:��_ĉy��Y���}�̄��s��pm�<i:3��%`�\.Z��e�us&엔����W��f�C��
�9�����H( ��1Fϣ� $W��9y!S8�o�����/�!D��?] Z%���Ș~�]�U��R��,΀�3�I�� 𥼋;��#�C(d���c4M��9q�ÂLr^ګf�z 1Gl��4,�@��;]t��MZfLm�=��,���^��?�7B_#Ɠ���`0 "K�0fî_�ߌ<�������J���[r��] ���Vŋ����.��f��T>�0c�����^�+�G<����-k�yZ�H�e�L�M�,������+U�����N7�\"S̰����H9�M��iI��m>s7Q^5d�s�&�x @E�rB̌NЊ�gR�=�Д�q�c=iqV�|�0��Ѫ�7�ߥk^�ޢ��k��������õ�M5����'�:��=�3��E�	T���M+*�� L����t8�k%<s̝п�9����@��E��5�!�V@#�c�:����R������j��Y�Qc~�*�o	�{I7u����L	�!Sc�>4�v|��ɦ��1���!)��"� 
��O�Pf�a��2.�Ĵ�}W��_�M =|�~d �Ů�I���)�����-P����R�y��Xӳ��L�	�}��?7��N����a�(^X�Jr�BG�F۹�c�Qe��8AL��X�-H�e���ay�b��d�>�r�[׉̻�9(�!�t���.��u�V�c���,v�è1h��˱w]C��=U�i�{��V�wJ`6H:��HEJB$8�[�i��+Ѓ�TdCƞ�b���<�U���c���ٜ����wR4¬���_֙*�u�����ZB�i���T���ߎ��8":{������2s�3�-�	λ�yI!���BX��4���9�!��L�rN鞳���u�[QG��l�$�H�Y��#��\�y3>�Gw�-ŀa\�����F@ �e	'ˈCg,���TmZ8�E�`�H�;�	0��K_w���9���J`�+�e@.@�T�W��ڠ.p�A�+�C��a,I��i`zȴ�)�2�����c�:vqbÍ�VPoė)�E?hi�I�!�>��4�l>���:Q�a���6��-�e�`��ի|��r�O�,!�O�u{=Q�!���`f�n��>�7��B�;93�ܒwG��[�]n��E�;c���L���l�Bz���v]��/+�C_�[�]��l��U���r�[�d_I23�jYz�J���ܫ�m@�3s0@ey��, �v�-�o ����1��
�L�Z% N�MȀ�)��
OM(4G��s�@��v������ğV���/�ri�hN6g_�_�ʴ����+��k(˘��������]k�R]_S�i�Hy������0S��$��星a{�xE�ȥ_��1��U�6-/�ds���#x��<,�a�����P}���ڒ �5�#QB�l�]EQ�铛�X�Aa�L�4A�Fz��."����P�H��fwj��@N�&1�����7`1�U�r��t9�w�ˈ'W�'�_�[X0#u$�D���9u�5o-6�A��P��@�u�J�4Q���c�# i���e��K�TA��E.��wH>������h$H�Ժ���������΄@�|�[��1�2��S�\I(
��8}q�A�6��L�E��݀���=ߢݏ4��?�i��N;fn��x�,n�d�%b�.���q���aPE�u��=�����rT�):��g�Srd���/����<�����
�� N���p�:��&��@��W.%��"���ѡ"�Y t��̭%���@|���}kv���5���c�Y��󍏌�+� ��g#�cF�Y��.�H��P��³	XTVG_��?�nV�>a�E[�j
�%��*�羀y3��_�6��mC��\�7�E�w�5�Ej�N�3-��8ރ����<����������D�yOy�i�R����~@�
��h�nLDKt�W��
%�Pƴ�Y&	��?�q�.��(�\���Ml1��I�#M�Ĥ��:8�B_O�d0�V]T`�ҥv`���O��ef��&�����W�=7��(�TB?K���7���8g����w�A��<��GSĆ�v�F��Nّ��J�U�i��{�Dh��纙ܓ�i!�Ғ��� �?�t�)!K�L��
*���������٫�KU�x+�@�H��b����`C��B�ݧ�ְe�(l��wi�k�<�@�K??��@��@��!���	أ�0@E�~Nk�C�칧-�#SCo��e#��q�_��qCt�!刽7�7��b��܏,�\�=�*o�7fC��Ǯ��Tn���Nn�%~j���S������˧Zw�������*�L�e���m ���Iۢ�m�G��w��!��aI��|�^�;ci������V�6H=�3���7�?���c��-38��hFzt�%�<��$\��u@{l#��K�2�|Y�|غGQ<E�#j\:O�ω�x=/��?F�D�v���s�ƼQ�P��+��e"a��}Fr�H��`�����o�{��93ÿk�i���&��r�A���g�;�]���Z5��#�o�b�Q�<�����.�1�����R(���%Z_%����Dx2<`.�����S&T)2��|������v����vZ2	�$ͺw�kō'�}���捡jp�?ջj-���#cy�X��`&�b��oxכǸ� �G�M�����ă�>�"�VeEG�	�O1?�K����uʬ��7��S�N���%��MM���D� 0e@pt_�鄹�&V�_՜@=A�����&�b�#��?w�c�A�+���<z�Q]���f��U@�W@:���X��2]��ޖ��Z8+�k���JyrC�"��2��?-6m�p3PB�k�.>h��@Yo�\,[�4��#�����R���_��C��U���0I���xA�j�	3��>e\�8<[�Ө�d����n|q��r�Aͨ�.Z��ǧT�2��
���As.�]jSfP���T�E�X�.~�����O����c�I��v���RV�pE�B����G��o��8�Ы!���t�]�E��0N�}��S2��D�*�ww�3�~�i�V�ac�g�~ �6{3.J-	�w�HW�ߨ���<���	Ae�&���ܮrO��ᩞ^�,J&Vt���E�y�e�{H;�*~u�87;|���۲���w	{6�>�jl��uUf���9a$Ya���[��f���wsi�T�w��ո]�2&�Ey>�.�i���w�\� u@�u��N�跐��yj3�o�£�7�s� e��U���&�j���27�y�&�=�"�QL`�ni�2@28�8��s�-�Bj.Nn:��-B�c�h�Ȋ�i����@"�X���.�FD��# ��1���R���~X5AID5]�n�K���`�����QƇ!P#3܆�X����R�2��a�(7��m�2V���fg6�+���c�A0+�֞䶤�PR���vI<�G�4�������a�vDk~�Id���r+�r +���řv-ӕ�K����׬H&��+�|�&��8	�%��z	��Ee:�]g�i�tK4��4����<�71�;IU��)-́J��/�	��яx{�̮�F^M�}���+�zD��#�ԣyd許�F��W|ȉ�����i���^�P+� ��m�bG.��Y(Zo�QS����ܢ��9��OE�rH��o��A	^�ի�Ӳ�bY�y�<�uv�6ͱ]5yrhW���j`�n��lb���$����3� $���%��oUyF��Q�� 
�F_ܐ�J�{�3�1�c�N�|�� � ib��+�C?]W��»�O�G(�ꥶ��j��ɾ�ЀCu�sk��={���B�"��TuE֊��C�a�wMdw8:�J�W���X�B��$`�hy�U�Z�bD��0�4焾���O�\i��X�[:ѭ����>uf�H���C���(Ж�L���>�/�Й�ͽ'RG�;w�nU��UL.��ku��`�J�1�f�Ұ0�t�8(��f�&<'* ��#O�	�Xq�L�Cc�^�'�~v�	P�x�&o����Ƈ3[��>��H����)�/}�58ߝ=����l���I5g�"(aS���k�#�郴��8�E�K�zh7�B7��P�oi�)*�!�J����Й:S�mӞ��p�{u?��3᤿*�5�]�ߖRÔ=����6|!��Q|��<l��􋎪/
� �^�˥B�ڶ��	c�g� �wLT�;Z�ů[A>�I�8��J��a�ז�T��VI�טR� �<�V?AJx-^Z��T����o�	���c�1-+躼ʰ(2|�5��V��Dڐ����V$��>H��8��#N���;҄u~��E��}�����>Z?�g����x"s�!×�c;���x�3�_ ��m��C����
��Z����t��PN�ϋ�����)!ӷ�;};ay�1�M|wZ�q�@�\�v�jVH�W��f�
�Л%�s>�G��;�j.�@u&���a�#�:�K#&�f�hƘ�W;�8��;��BBl M�}�H��=:ؕ��h2$�((��A�-�9n�.�C�)�o��U�@��u ��l#�B).F��!��Y�� ~��(�|/,HNd	� qT�0�'���F"��M��@Z��Q�0D�-w���%D6̇��D�u�\��<���v�pkY=�[^o#U�j,]H�=fs�Xh6���F�6��g���B�3P�X��@�ϻQ&�;ۭ���dV���I��)�f���"3�^dbZ�h�n�S!U`���8�a�����;�BH����O��e��j�U�h8�=�^#�J{_e�������-歰�s�J�l��2:�2W�G�O�f�?C_~�d��l�W��L	Z�#�����/L��G����BF�ڿ|���	#ȟw�/�e�ӤS� �M@�w`#s���ײ�nX����Q�D�\q��M����M�*�ʴ-��`�/�wӚ��e<�,3�Uw�C&�G	ܿF �ق�}q\�%��vPzq��w�C�+/�׮>�4>��m$t˳���C�3+�yZ���T�!͹����\d�w��x��n�9�Ԡ5�L��!.\�BH*�e9�sgTYL%�)�|R?�q�Ȕ���/��qބ���&�E{�b��,���K�.Z'q�(�Դ��T�ߚof~�aˑS8ƹ0PW�2v�����3 �S�mt��}��ݩ���]@Ĥ7�
R/�����l�T�:5���=�V̢�F8�ɪǧ[�x��ϴ;
���lL���D�xN����ϡшK��r���O�->�odFːQ�-� PF�K�<��\��{��}�ޤy	~��Z����יY*��E��a.�vr�q�ek�Ԟ��BE
��4r㺯O��!ǻV��N,� D�U���#������b���?�����\*�U�D)˪>�I�!eob:���Y���g�O� 7P�P��1���r���x"j_�@㿫j��޵��+�?��E�k�����JG�~>�[^y�b�,�W�N'�a,t
꼭P%�D���um湳������ F�@��*��1����X�`4;�l3�\��v��� ����$��ݴ0ЛDk��n�JS�p=��e�2[�&Ɍo���6�N2�(y�M�!��_�����]�������)�������M�ߟa_�tEN��X�N�Z�L�zjp���m�'��&f���JEj|y�<y�:�Z�`��t%N .���.h߁V�0��F��)_�-h��d��cR�R'�S�
� �#��'T��rE�A��յY�MҸ�������~��x5���� �/_qq e�I�zp"�4�7$�&�j;�������p{��c7+俣'=g[��-\�U<���
�e��h����'SB�*�4�q�NtuC|M�OHi�|��s��d��~�����1��|� ��/f�#��oX`�;�x^�&V]ó���=)�2�а3ۧ�L���T�z��/�Ŕ�������������0��M0�����_�����,}B�R�gJ�ˆ}-RG3��X�P���YJ��Q�%��R��M�!ޕE�j�� J(�_}�����= _���3��$�3���m$$:2���A��W��ˡ-��!(��W��PFI��v:�JS�-�.�k�L�I�ׄ�CO�����·!��9�5�7To���nP�j{�w(�tĴ�)V���������	�x�@J��]��*�z��CV�dy�T�>�1�jx���c�w|K�g6K�f'<_���ٯ�
���ֵ��g�i�D�p�"�'�kdE�O�u���S�摯Q{D�4���K޻QRi�6`6�u�d�OMo%�� End�Ay� g,X���>F*ӌ4P��0,�H�Z ��`D,j�l��A��������g�����#�^H���;N~X���}��Ac�|�~��sݒ����5�#<��|_U���TXc�5�ۃ�{1<]~�"4(\�u��z_yd��G��[ YPؾ�� �kj�i�z	���V���͹���C��'H6����\����F;!��(�g�(��dȌ/�d��v��oІ�,�!)^��3����Q�s0���m=�^nb(QJ(Wh�9%gu]������R��wmuځ��.�Sd7�SB��?X6#�Bd F�*��`�Z<�>f�{�xV�XsK 3�)S���FmQ�����ݜ%4�Ź����x5�?{"�o��tG2Z�S���%&E���9Q{)�Q���,��؍-�3�T��T�C�t�EqP�*��x���*���n>9�.�r��i4��AB��Ypt��c��m����|˶�T9��s�Z8����n�z�H%�0����;[ڙ� T	I'���L�	�w@l�Sj�kl�� og 9����\9�Z3��ێ2������@	��� D�Jh%�1�t��D�ׯ�m2�*����i :�)o��iC��p��0>�<|���0��Kn/�)��i|��<�k�GF��MZB9͔�q��!������A�L`|i��<���2����P�!Q��*#a���y�/x8��uJM�)�!���w�g�`3j!�mdN�zw������ՙ�z3�5fS�A��^^D�dxr2��Q]:�&���l�+�@v��i�!9< RZ�&(���\�a�S <����М��%�J�<��CI��u����]�_�C�B�i�1|��Z��x������z��s$S;N�v��"��w�������H�R6�ꧬs�ŏm���<���V{EF���7�>I��{�Y���#�1�T��0�+M�C���&(����nEL���.<{� \u�@e�����W���OT�n��L*���,b�i�F�6C?�g��O�^��+`��7C;#��:a���ɟ���=��	�چ^���W�תڋ�dJ���#.��0^yJUF�XIFFJP+{mh���F����'�|�ƥs��D��W��Q�D�얗?�#���Z�'EMG������O�p
?*=�P�t��������lz��gu�������q�<�� @qe����̄3}�e��j� UK4��D?�0�0������e5��ˊ�t	e�Y��T>���V����.�]j���-���i��d��!6,�~t�9Ƞ�+E�s",�����')���WvB�h�����:�3`���K+;�2"""��ﱸ�Zr�3�}膄H�	+:����f�5!�E�H�f���,eP'*7`>�	S�8��Y�On�͔��x�ҏp��2��O�}����(����Kճirٺ��ֲ�:S��W�Tj�Ǯp1�� ��UI�Dr��]Rb6��f���K����IӠY�KLR�5`�+�9�m�O:��͓i�@��_�0ګ�����m���QB���.!�u��2����}'n�^:,����;u.h�5�;�n��=�do��Py#����F���{&r3C��� ��1�x0�_�1�g�`�nmK���o�s A���P��kWp&%sV�Ke��Vl~:�~6&��8_��Ñ����o�[��kH>����A;��$�hx%��6{.tO,[q��n	�F�6���q��nM
�]���ӽ�ՁWu>׆C��iu;���ק��ML����kA���=�D���'�/pJ�l�s�]꩔DZ_��o?�*{�����[�Ŗ4[�c�K�4D'L?1&� ���՚¬CQ��ۉ�A)`L����5����3M���Gw#��X�'��w��FR2Z��i]���̀裦v��9�9�����I�}�*P?�5�;���>q��s2K����3���]�W�_|o������Ї�ox�Y�A�FxT����S�P�+��,�ª,�b�sι�k���[�)��KH��q�������~��'�!N��G����+���6��kp��=�z�WO��$��' �l7��r.��!����6P�a<��|A�
���
�v˧��"P�ܫJ�b-�;����f�n�2��
Gj�Q�zmv#�rn=wZ���e�}9�����A��8�?j�5F�\J��x�`�L;����`��S���3��
����v<8�,t�8BT/|� 01&�c+�P�d���Oy��R4���_cdZ4�����E颃��G��~�W|v>�H�2+�e��b�\��B�Ȋ~/�x��#�RJ�B%�צ��ٞ$K%̔��Ql֙���©F#��pd>rA��n��G��%{�����~2=]�N��Fg�X^J.y�u�8#����N`� �W�荬�Y���U���/��:fL�b����
Y;Z�3&a���]W�@���p�cͅXcM��b�Uf������f�z�>�i���K�S�w7tm+����*�.P=F�Y�������0��$�T�j�z���(g��Ý�	9���,M=H	a�_�l��m�R±�2h
a�Z�HhD|�b;���ϔ��$D}bA7E�W�U�B��N0��ĳ���ۗ �SP�ѹ�ez�;�6¬�x"#�$G~�����@��Q��-wy�XК�$��*�ڸf��=?�z�	,̻݃����H�"ZX����)����c��)�Fv�2؀o�Z&��wЗm�J�9�s[���B7����h��Њq#4�r9j6����(�� ��h�S|��ox��DO��J�]"Ou~�]%��1�+Y�J~ �����B���D�)�5"�0�
�'�CH�dw� +�<���JO�2�7���$�����("����	�B�Ł�Urƽ�c��<��X��<H^�ky�9�;����lІ5!����z!T����ם��bC�N�?��c_t��ҭ��R�R�~ ���.d�}v0Xf���0��	 ���e��8Z�O��t�׾)�`��n<��u?��$���;�G�2��ճ���K�=z[$��S8�To��`�')t�c��k��G�L�:�@5�d�ܛ0��������?.��ݾԴ�I+�*E�f���>�`k�lq��ք9����^���[��ҥ3MG,E_SMQ�.PxN������[Z,�vx$r�ݺ*��f>J���;6)LV�m;(:	W7"a�ܜƷ�J��ٴP�]V���V�1��M�۷0���)	�]8�T�^�xT
e�i��M���܅�
���2i��D��� ��\���&ʿ��\L�Z=`���M���a��������b��뻪��G�$g�n���PB*ᐾ�����R�>���i۔���"m�c_��k���z�G�hU�!Es�Fm���i��mQ�M�zv�\���T��!��z����9���� ;+�1�* ʭ��A����*�x1|-Ŋz�Bn�en�o�LI���}F��ĬJ�5�>�8 \}GK�yI@|�x2�a�MX�$�L���1�	�eR�Yj�F�Hp�c)p�o��\G�$��_� Y��,�%7��f�y�w"�j� ��i�k3���w��#�ծPI��7ر���L�B�r(�Y����X�� o6�7���L"�u0��0���>+_z�y��ŢK�Ã��@	m�;	�9��<�*l�"A��*��,,����Za�:*I�9էy�����g���6��X������v��2��N��`���f��	�5��Yg*:�߁`�\�@�.a[1�������da�󰙕��;�&<�J�Mi���g���r�0�0\Ct�v<4����PZe�>`�-��A�OE��
G�5J�Ϭڤ�tƔf�+Ч��Rc���'D�F+�(��nyte�& ��'��E��٫
@%�.'���V���"u�|xV�� ��钫o�gGѫ������%���gv���*�b�:��]`c d嫵+���T�3v^�������ȩ�j臑}��S��Zg�0.U�3��2���(�Kɞ�~,~������?^3� T�]���ಯ��L�d4�]�3<�6�.��	v��<s̩F\ٌϊ%�xCK���H�.�)���ȿ���a'ma����~i�D2�iy�Q3%��̗����f�����dI���8/0?ߵg��$�]ĭ9H V�Q��b{�OZvVo�g�5 �k�����;ص絯��5���<o�Rg����}� p��E�_#v�0����� �s���2�k)-Wo*p��O4�t%[����ۚ	U\洁k�-��?��T�P�C�'�X)"D���|L��/���!P>�<eE�|��1�eC�K��Ɏ%���A����(���+kI�r�ǭ�/���w����jŋe�q�/#���whQ��L���}�N�{T�J�h���nhsM���4{��t�j>;Ã��D��`Q�4A�fkX|��Rz��&�^�R����wp�n������ъ�+��-���;\�|��#�{S�f�0P�L���Do6U�C�%�:B*�?C2�d4����F  �2z�ꢀ����mمN�Y:�Mw���!m<�����J��h� �a�h��!�(��O�r݇�'�>���T��p�"�e��|�|�ܧ{�;ǂ���$4�CW
w��%�F}����'�)�J�E���!f�H��rh'��^�Q,Mޖv`��o��Ԝ�eq��~�fsZƆ�|2�c����}薵�85���kk���/2t2����E��K����t���16v�ྵX�4K=^m��k��[j#��ZV�,�ʻ�
��jmd�{cݲ�n������������hy���msu�Fd
yI�a�澘(��{�[W�q?o�"�B��cI���'D�Aç5F"U�q���ˉ}:~�l/��x��Լ~,�����+!��=�G%��+I/�l]�������L�Qˊ�Guuz�9}p?�HG�zB�73i���)_mW{J�ܢ;^V��5AyE�9��	k�׹���2nV��qgHȏ`��MTvA�Ž����(&X-v\�nN��^li����D��Җ���VI���*�?|ފ�&d#j����Τ�0VSC�!���	p{��g���N $!�*���!�S�i�9n�]��q|'�ʨ�j3�I#��-è�|�����d9�u��a���V\���N�]� |^�~������/�	}eA�[B?���A���]�Z�:�Ү�>�<��⥪Tj|�d|rt�Cl��jG���B5�,0�\\��2ŎJ�ד���<ѥL� ��xvt����92�n����ۡ/�~u��w��ל��B����i����}������p���C�F�����t�[|&�#A�㠞�Ҕ�9��!@�_Y�ѡ���U�aL�m��@���<�uC~M��������G�\�E�^B��w'�n������j{����GY̖��@0RcF_�j�w_���|�`����H�o|�Aƍ�%�z�q/�>T�ܵ0v�M4��$d�;��0�[�����:�sֵ�ѥؑd5<9B�h�_��S�\K�Es�$����X���WIJ�r��؏k��v�����L0�N˺�RQ7���"?~���a\?7܉ڦ�?W��|)���6�D�'�(c��hip���;��
���mP<I��-�FG�8� f�������^��ZՓ���W^ef�F�O��d��2��Vn�3h:� �yE�k��S�L˕_���v�$Z���m��[����&c��7^Nc��6Ơ��A�xyM�x1�����]L�z�pg׷}+m�h�y�P~�{���P��k�H�@|�^+��L�x�+�f�e��.
�M�G0BU�`�հ�y�@X�J�_�v�W�l�ktc��`�-%K��!�|bt��@�rω���o�^�B�8���`��R���Ʌ�b09C�_Z�bE5,$��:/Ш�����鐽�8I���޾
��Cc����)m�}A�%�w<���נ��4�(�0���G�%���O��?��r$k�J3�*��Y���Nڮ���"�x�Jo�dp2|6I�%�)�LY�k��#���ѽ%���g��xJ���E�C�/���8-ͩu���c�K�X�;����/���$�SQyj�%&�jKC����W�5�<��k�������Hf�:�� ���.�£c��m���.O��1Z����(7+w.`��mT2�)�'��H\��q�N((�% ���?d��j��w��FX�6���?g)t�#@*#��]9$���o��A���!�b3~���Z����Ȋ��Y@����'�E�Un���`���9�uFw�OxN|�]dŬ�|�ϋ�Y���c�&6�f��G����e�Q*���꿎z����C��j�B�6#��#
C�[`����2S���"��"�$'7j���jԁ����/�6�U�\��YE��^��B*�"�J	�Pb6i|)
!��di���(G[i�MB����?�W������P��tV������D+Z���/���i؈�Zz�m���gO����b��^����_�8,iY�N�_�} �wQ��ی��Cg̓x����ʣ����1�߂�e��JX`���
\��ñ4���_Q�%�I��p��orʡ�D'E��z�g��7uK	�Yz�����s"��Z q���� a:������)������x�����=�s+�!�N�K�\#�p�d1����+F���"�H���%��];)�2/��~ߑ
\\`��F��xj��������(B	D�%��_����'W�.i<���Ų�2#�h\��d;�_grں_"5�LL�C��D�kn���8�t��G�I�������r� q/~R��R�2��?1}�m�>����x%�cep�B�YC�:��|�`"���S$"?*B�]���K�B`�lU�{I�m���*�K$�|�B@�/Y]dS�a�ۅ� %���1�7����S��m��E�?S��y�S�(��v|�����U4ji��	�+%q&��WT���$8�x|���$��)&U�4��(�7A�F���@��C�dͮ�����?�ؖ�8��
!�v9�~t .�"�z���z�͠C���eݫO��
m��+�V��
ƛ8����JhW�?(�a�U��.Vo�/�n���Ҽ�i�\��;�1[��l�w�>Zb��Vp[��9���Q?Fr���%8Y8ܦF��}��TS��v�v^CBJo�;�+�ck�6~�,�H$0w�@��bh�t�W@�k���y��策]ό��-���q��`�v�]���b�)h�Ռf�ON\�xZ�!q��̿R{����}�$맄қ�6��<,���xag�<�;�����QU׺�{w�in� Q�u��`�'�P�ܝ )�8����	Cp��!�V�46#��B���V�+I�g\�~�$����q��ڎO@�78C����Iy�OqA�4J�՚ME@���~���qZYp�BëC	���#D؇�ˡ8Jq������]���7G$4�N�UAgr������i@��p(�3G�����Z3'Y4�:G����RYpYc��7ǀi�l�q�0����U���)kE:�c[0ŵU��v�� 3��L]f�"���_�:`u�nL�qV;����2��p�
=�-4o�x�A����c]�?�8�L��k�z	.���U�dVI�괚v�`d��'��?�!��q�F��Ɓ+؆l��K�`y'�5!%����O�y�^�Mz-SfG��EH<נ��Qf�#�_��ИX&*7D�ܜ��П�}�x_<n��+ZL:�_jf���P����*�V������&�}�8��.3`7�RT�a�L�Ti��h��ZU�;�q�g^��ȍ�^Z����:�ɏ�ޅ��
�X��B	���g:�!��R�wև� ����ſ��F�A&��?z��nY��z��P���[��iW�.X�u �YBφ3S��(>EnH��V�e�0��c/h0��-�	B�'�Gyך�S\C��yi�i�Kuqt�z��j��
�K���R�����&�r��E�@���%��DN�c��OR"�v �F�-�-�/���ܞ�#��ҝ��	Ed0xe��h3?�v�/�r
�Rb��}6�/�r����yx2�,�~Km���[�����A�|���p���8��}7iI
�N�±�`�^�����@��gS� ��+�2���'z�Z�O�|�*BK���Uvi�,���P �c�&�Ŏ�U ��I�!r�9Y�2_Y�0ߋ��[���O�Ba^�':������O���p]L���k
��E*V�u�z�^�7��3�����9&�3PV^�A�@5���K}P4�3%�oa�����fP�3׉�0�_W�v-ۊ��t��j�@ �o@���\~<+n$��j��C������|M����Y�����0�.�z3��]H����>_�N��{�BN	Ѳ{��(�Q;��_
�D��g>�qo�A�-q��2�Y+~e<,���b��R�wƀ�:���آ M�qB�o
!�[7��+뱕L��$\�
d��DU��H���?�>LL��U7�`MC C+��2"Dv���1K��mߧE/��X�Z�6�p:�mR�9�0)O��e�/�?����T�x߫`2�jHZ�e=�E K�l;z��PA�8�?��-��nO����
�m�#Z��8�4�a�@�~$��p��(6�X���>�qc�z�r?���| ��.�Ɂ��|�;��O�A������I(<���j�*�=q���g���_����l��Qh�߉	n�X�t1g~=#L�'�}���5��ڄ��j��'��MeC̋�[��"�Q����[��
]To0�b��2b ��Bb����6uC�+�-�/� %g�X��4�f^f����������%���^Z�[�k��f��&�����}���Ώ?���x�5��S��̈���Dwc��{L�����Q���Ӊ���nr��Ӊ�6˹��
H֋�UK~_�)��c��X#̾�'di��G��zC$\�nL��uf��Li@�Ŋ;���-r�������A��$|wgj��l����EHOX�
-{ ��Ѣ�.����D�k.1���"�!�I} a'�klG��}��&%���>x����3ZҀ��I���_,�o��ݖ;A h��Cc��w�#9{����5���e[)�1��,Ę�_�u���Ӌ��>Ӫ ��h�O��x��>��{�,mP��9y=<](�5{��-y��}�*�4����E�Ϛ��m�q����Q�iRΠ8�)�D�V&�%���^�tAU���R��T�/�O��=��p|�0��$���=Z�̵:6�Ipkr��O�F�WZ	�����wcـe��JN鼬臭�_�l����3u{�(8ӏ*#.�U90Oz�/$�w�ř�eI��n�,��q���5��$��I���
�b{���.���k��R/��z`R�Wt�v4���𡾶�8��{B �u>��B� �5��C�z��&�=v�?t�f<CD"�5!%>�/WYp��p���(��ĳz���Ժj��+ĳsɖ�e
p�W����fe�g]�nPsϭ�L�n���:�C��<����x[9�pВ����	uo��;��.�"�\ w�7?��]�虊.U����J�%o�t~+�>���������erd�õ�b��aI|�q,n̹VS��������"g�������e9��ъ�xo΄���a��R�
��b;p�߮����I}^P.����d֨���޽dw5� ��5dja���6=��ʾ~ip���D�b`��1�������.H�����֟ap>�~2��[�쟲x?��a���t���>�=<i9�ÊՠϷ_U�r���۫�Ɏ��PT?h����|v����`j[�aR�s�7r~��f�J2pa��[����z(r#��<����l����4V}̓��c���ز�^���#�=�O�d�-i�̡kQ��[E2���4�E������q6sW��.�u�������I�-�@|�e����ឃ�f,�6�o��W���f�X�0f���<���X?�AqW�!�Qyr�s���O95���-j�p�I�;X�����}2�~�W6�R��^B�qx28��]��^.$S���UZ@�R8Q����2��3�� F76X2�g�a6��N�c��`���M��(,�[�X�V��e����~����V0��o�����H)��O45GN�S H����lht`�����eL4s޻��!�@V�o�%�trj$�,�hb��oC���Xi��������f5��#�����MtB܃y�aH!
L)X�
K>������>��Yjp�pO�!����x�^�v}I\������V+<ʈl���#��S�<���������$�!�_�BUm�=��ޯ����)��_W�\q��c+���`�6;���g^�oT>�oM��;x���J[��dV��3�ƞ�Zy[�_�)c5�_O��YD���K��-��_#�����]��aU!Y`�63$Jf��&�wgw\\�:2����[[k|K�ZF9��d����2�ڏ���eA���h>�Tp	S�RĶ3�T�6�Ql3�\�s��m�;�+��+ř ��Cur�]�.f'[X{��g[.�a'g�
���9�����a��J��@F�\�Ɓ��wBDNS�BH��7In����7���ǝ�RC�hJ�\X� �b�ehq���=,"��T�:�B�N��u��L@�h���0(�ҩ�iF�G�C����>ǣ� j��^�����E�aV�����\����j�������61ɡ�����k����*��#�R��yXIi2�Hv���%�:�X��!Y��Jz��|�����Z��$��ma_u6ˠ���ay�P���	�7U.��ʬaUf�E�*B0�/�>�����x���7+�,P�Ou)u�P�����-5@
�#�3ٺ&��y�#�x1~�ڵ6��g	��썑_#=ꪢ�q�:���҃9X�:�V�~���q�cWɡ���8)�~T�{�;9���%�6L܁������f8j9���a�*��=t[?��������q8�Ų8R���8����r1W�X��0~�n:��NKCN�u�w$~z�%�d���U,�X�T��ؠ q� �lGLo�qw���Կ����r: -{�SX�햖{���x��BT5�T/���!N�.�����1h%��hT�~�6{r����u�W=
j����4$�4�KEq��Vڟͅ��|��zb������]�#��GJ�z�__<AV��~I�^�:완i?+?^�'r�.�K6໇B M�Qm�y'�z�_g8�XF	&wۆE/�˓��\���v�4��q�
�<��8@B*A�b�ʵ���S���iE�%�֬݄r�k�!�ǉ����OM�9�{f���6?L����D��LGt��v�\�<�<�Ipw�b�c/-���FR 0v3��������
<�.��H5�.���:w�S�sQwSA�:n-L]SD�S�4<i{ �/�󺰻/f,�*:�&˻�J,,�ѻC��S��ppS����}�; Qe�#��}�t?�!V4@�<���A�s/��6�v���{����1q)�PH���C���:r)z>��]�6:t��Q��������֭]����R��:��O:��c���i���sQ��L����p��
lNȅSI��l���_|��])��(V�I����z��&Ծ���S	�����E�!�;�5><���j�ɢ��5�v����O��
����Ș>e�I�������.a�S����gD��~ͫ���J� @X��KC"���{�f���aً-a�ߑl���DP"sE[�.��ʵ�!���^C{�"F��6|#mmH��S���i���I+�М���,�o|��W�7!%"��\'f���qE|dhx��x5���G�\1 �x~�V0�>G�0�r����4X����h���O���7��K�g�vg��!�Lz��qOX@�;�un��4"���HB�[��ܐ���K�0V,�!݋^�[|����_��Ħr�졮��`�]�\���M�f����6y1X�^'B�(��7k�X5_��u,��~G��k���=�DQ�ؤa$���Q8HC�h�h�.��S�K{����@hS2�C�C_R��|r�Z`
�mb5��T�S���򶹎t	�'��*4��������<lx�ǁ2Oh��Cڔ�����7���Cു��:n�ź��,7QX�H�@5�02}���w���\C�m"� �)�]Z�Q�*��Ty�������Z�Z�J�5�$+i���cc*��X��d��i�nXY G�lT��rW���x�ʄ��M��d/0Ϭ��Y�g9��1��
2�9��.�|����C��2��uKB�;L� �GZ�1� +�A�T����0Jf�g\L�	��0^V���V*rY8�H�nD[q,mk0t�9�\��c�h�Z�E����񍾶S�6Hb����v@V����=�FQ]
8��N��&U�4V A�`�ʌ��;�!Q���+P�J�5R�(�j���O��������)cg��ʋ��_3���7��!}G�	�Q��ۂ�X�����*?!(Z�0���,�T+/��^`��+<5������Dխ&�	��U�"��La#�\%W��{R��m�ݵݞ[���]���R�J����}�2h�����*C�+Ŕ���ȍ��I7�MF�c�"�!斪}� ,{�{��!���`���j�!y������U�5� 3��t�5�I�}��U��y�j�- M�ʜ%�`�������m��9dl��A0���ӝj�W@�[��GcE[6���X���O�}�# ��ʖ�l��\��l��b�T!� ���R�B�{mLGM���h�ai�"x\	�yX����G�����ɐ8�-���x�K{�q�^�-����4�@R���9}��`ш��,��3X���ؘ��[�"��������N�c۱��	�<&]��U�x-����c�P��cr욙ްF�`���D��3˱#qѰ���Xb��8��4�ק��޶�;*F�w�X��d�`���hol��Z��6Q$�r���J����F�B�*����3������P���䂞Z��Ȫ�����cs�S��v�>�ާς�_���[n7Y�ψ�'j=�do���3�]��z̀�;U�5��J�v�,ɂ��[�:M�wC�E��+�c�y��̙o���1�cF\����9Y���2.NO��/Uu��
{G�H�}x�D�����n��_L���E�&,�)�PG�1���8�����NU�\�c&]O+I��� t��&T���%�{��ЖcE?�MQ��4ɸ]�ﯪ�MS�Ԧ�D��	D��y^�w]:r��t2]�����WR�/�V��_h|hz�я�I�)���B1���'u��(�H�<g �vL~�El�g�&[��`�Z
e��X9��J����1v���������Q⃄�#�q���y`&�x��VUs�}&$*��a\G����,8��;���\�̓��m���<��_�oL9�bFjaWM,��s�O�V�y\IxBV�	�bau�@'�w�k�9���p��&�m����Կ�E��G3Ɇ�P�rt�nMG�j|�TE��A������}Q��Ƀ���@��(��8���L�%á��c�z5*\_w�=4����*�C�u��G�G %�g8n1�;taFj�e�=>��n�/@��%0`e*v/�j#~��p���ʸ�[�ݣ�n�'|�g$#&+����&r�Yk�\����Η��	�/��U�hօ�<�뵁[~�Fw�E�Ĝ���#��_�0�-Ĝa�M��w�����p���4�i*�`d�U��$��x��41���u%�S�Y2v��;�N8u醥0 ԥ;@E昕$_��6G!8�����2�����A�2
��Db�[)�-�kr+(���]���U����Zi�U�]p��H�'xzʥ+��u�N[�e��8��*G�}�@SN¦����+��P�d�qk��~�Q<��}���S��S�2����ܪ���:����~�y��3�Q��6�r���OmEh�/�#� �W��)"ŀ��Ю����c�DB�����Q����v���� >E��,RNTZ"#p�`�kޘ+d�	\4<"�v���8܍�8����9潖�e��^!M�tvR#�Ss�:�Xsl]�����r��v�m2��a�}I���S⁄��]�����Z��5T6�2��f؋5�&.5�~��O��C�;޶��̰`��\ۘ/@O��+�E`�#W�t�s�a<i~��*f\���L���*O���
�fuq�/cC=�&�S34v lqt��N�<���~�j�m%�X�1+�@�ؤ=M'(��_R���һX���{�����:�ۅ���^'��"���9;�_Y�_s���1Ҽ�uhH��u��Z$�g��@C��8�d��|��E��
h�
Ө�F/0"wZ$cO[�Y7]A�M>�k��v*-Rf��<���M�����6���}Ve��a��C�WN�$|�H2���� ���U�U��8�/Z�u�Rn�;���E����q��V�Ao��<��{	���S v��,}���GQ��Pϧ�$B��W�jr[������{@�ZK�q��q���h[-�"z��}�B_�l#�@]�#��葀~�!��7�z4�9+^
�Ϳ=P����Q*���K좚�U��4K��&v{�c�ڸԽ���X��j������E���C5�1��4~�!��ʭ�-�B��L$�}�T!i�Z9��F���n�.��n7��%�E�KK�bo��Y�sxV��Ǒ��<��}�����9TXm�Kʢ�X*I<�R�daJ�,>��H?�f.+Z@���m��Y�=�Se��'>&g�5#�{�}K��+@
��� ��;����ů�9���L@$�E�W�W#�:ٺ��L��J�y���h���Ͽ�$~PC����S�J7���MfdMϵ����	G������&m}H��mߪ`'y���7Z���x\�`o�n�&��Cv:��˖> v�-��_g�@���B��(h�|H%�v��O�mɹ�o_�+خ��/L$J)]\���{���;��a\zގ�=a�ov�4�$q"�H/��2�J�Hbb�[h�E�i�����f�k�����E2��?�a�Ȓ6�CG_v����?E�$���J�J����������ιr��h��k� JB�@��!|=�#h�sg��`J�Z��Յ�f�VBND͵��]�"����t�2�ဠY�$�D��G�C'l�Ř)�M�a�!�
k����#* >�,�v�*<azN���qm��C�����.��[O�r+&��PD��r-6��a��r*���G{#O7u��7�?'�;N۾�?���#����wח0ԭv3��h�xԊr�\�#�O9@YJq2���Cu��N��	���>@69���
�9���F�LN���0�6V9�;:���#T���@���֪��i�f��t�Y�
Ց�%|�IM�|0��F=����Nv��9�؍E"�`p�2�%Dk��n}�Һu;�Y�"�[��ȌVq�i���ZNxVP;�Cm1��h��?@IK#��\����u�ٱ�ԹkI.Ʉ�J��q�>��|y�q25�롓�L[0hji�sfn=zYw(���&����� i��cD��k�ߣq�)�x]6�w��?9�O�ŊG������v�!R=�C��'_��=�u����_�{텥� ���/�k��8��4�Ж��D;|^�w��{�=R�����;F�0��V��1"ɂ>k��Ź���[M�%��l'��{ó^�᭔*�A`����5ϋ����<ư��-��2};�z��i����5�H[�'t�<pۣ_��m��"}��>���fi�t,_�{J���	�'�_�O�/K~0�Z�� 8�Mq�w"�,��}�+T<�����CźZߨ�C�F���15�2Pa%`"�8���%��R8u���R�����'oO�ܺpu��O0=p ���HN��.E��fE
MBʵd�=�E����(�B�bC�Ɠ�\o���#fa����յ:J�9;Ô��=�"�����n��)���eQ�9=bb�(���{�'o�i~3_i˅uD_`�������2Ckc��7��}�ӽ6_��+_���EE�};���(��A�.P�Ȕ�� 5T���t'Ǵù�U3��Bl�t�n8�1�n�&3�Ă�C-��F������5�V��8���u�����o{�\��T�	4��E���ylH�#��C�R��v�L`���9�[M䵖j_���RR-g�a��\��zR+�"���ǎψ�ʒ�Zk7�[�\�e���%�~�O��UΣd�n���rg������M������p�g���6�F��]�B8�b�<Խ�q������0�PF���S<J�!����o�F�&�8���oa�U��7�7���~��l�}��cTIb��sKG�C�<���%D�W�W��m2�p�)Kp�LV��+�Y%݃:.�#a�Q�t�5Yլ՚����kͲ��n)|b�3�ksP��}T�������lM-������e��U�w�R&�R�]~A��8t�{����4�;$�0�j���d��[ �q[A։���������}S�:VD����T<>��]��<9� o��}.;�1��`�q"�{M�*��ߘ.I�2�����>V�����|w�?�_|����~�#q�UTW��z,8�k@^�?	�5	�+����~�`�����"g�!!h9%w���sP���n�^zSA��>�����O��'�*�t0�ʼ�$��10}S	ػf�e6�v��NN~����I��EE�.�R�4���Y��	6�%z5U����(O,AXO#E���˝�@XX3�������c�ڲ^�yi�Ӡ�ranL�h-�*.��|�OR8(��<*�bE~�H�p���ÂDo���w�k�4�<(t��g<l�"�(�l�vMOʫBB��l�y\Am���'"M������+���ѪJ<�j�7�?� ��h%�Ze\;���#s��D�B��1�P�m���mB�M��[:��@:\��_���9-.˨�q���!w�/_��n�nK���_EhKWF>���Rc�OR���͢��7�֕�/2@�ʾa!w�	:��,I�����U���KV��C�.P�ϸ�.3���u����	�6ԇ�q�=J���Q?���/�k:X��gG��6Ĥ"��v�]���HW����YL�>*5kT�v5�
��� j��J�Ϊ���E?M�u��z��������n��8�Xi�~���i�B�(F�'`�ĦM�YA<�gv2��>���r\��R�I��k�Cb5���ʣ����q�J��A")�����bid$�&�_I[���~��ʲ���a�崨N1��-jy�U���SV�����ɞ��t�*�Z����C�l�S���4�E�~� mm��5� Zn*��=f�{���7P�M��Ǉ�&0SY�9ʪ���Z �n�*"6ü�Ȟ�vЖ��{����퉱䪨<w$�����8R��5)�2G����4E�K[x�a"&ɏh=9�]O�Ū��<�	_���_�p2Z?�O�!J�Y
v��P�P�����.��٦SiTn �'.n��Xo�o���^��������ҁpX��uZUw�,Ο+�fޢ���;�_7t�.�a�����\���gufHn!*!��z��<���d�����Y���n��k�=g��Q2mT�~Q��U��8�Y��"{�$.Y�v��!˛}/r�d��[o��4p}��Y).�U����:��71�sς~���)����j:��Z�}���]���B��
wio��G�p������$����R�R�Қ!��N�!:�;�|j��*{�L3`�^ի^��x���L������(s��Ü ���\����wF�}���c��P��5�s!�]���et7���ä���E��4����a�VQ�c�)�+{����Q�(�� \��D�_��~E6��L#+�H�r)%���L��OCwƎųr|��
:8��*+W��f�hm�S�Xj��F��\�fw���D�O|� -��[j���Ȳ�b�#���4�6t=y �����U��Pe�"s_��_Qq��0T,26�il㦧��L��	�Ά���3P��V:��v�׌1>�(�&4]��Y��J��Z�;�)=�&��Z��%e����{�x��ƥ�:*��� �E�a�yo�o&r�J�i5=SyN�m�3�i�~ʂ\�!�τY52Qc5c�pC����])_�]�g�LJ,7;�BX�����@����/F�p;#�����Æ���}?���Û�8�}f�P=�eB�ǎ�P
������B�u�-1����Ǿ���E&����0v�JzvW�|��.���D�A�������<�O<Yg��l��#��>���{��z�+X�<�t�v��$��
��,�L[T�::&2 ���PF�\�R�$L*}�U��˦�����$��W�����t�h\��u��Ȓy�X�݊�c�}T�7�F��'���XA�p��#�M<ip����Z��[�2���4���cB�"��÷=�#�:�~�R�7�C��Z0|֥f��%�<���7��g�;�x]�F�[g��
hX���ʩF�,賗B5�2q�;w�0:��;Qt�x�L�yPg����6_�a�?��c7pa�5����͵�%�#/���*��oH��}�}�� @�f��~]$3p�$����z����_�=�i_��6����G��-����)>p�'l	�y�?�@����٪�kT  cͨ�Mg����x���t�.�R1�(�A��HҊ+s�k�sr��!5��+'�V&�-��5>���>�>$�v7�a�sΉ�XDD.�:�	s��?r�kW�;U���k��X�Hj�,����<)]1neWB|U��lu�Ζ:�G!p����_�y�Rd}7�[�<p������bZCSU"@�j ���9<Z��E�dLV�"x�B���
v�SY��w%���񿳋4;���5�r�/!`d#5�y1�$�f�]XQ��#�?j��*��d^���Q�y~kF��6+�0�a�f
S�'���s�p>k�;l٩͜�s�t�r#�C5�0Fz�jw��x�J�V�~�v��MeCy�^yg���B5��r���`�׃��1w9��X�P<B�C3g,��}�L���X�B�t$J6���ȗ�d�H��b�4�<�����#So�rbE��w��g(�gV���ݯ~5�f��FJ������.5C���=ޒ�� PW�k`:T�	�[��D��h�3�Ǿv��X�S.�n�{Ȉ"^\�/0I�`�7�OWc�"���5�;�;e�Vp~j
䈃����'��G�M-��r8h����t��������%�����{(#���"�T C��|+n�([�F��S�w�X�Hߔ4өV�D�B��-��	߁E-��"/b�`h���X�V�_��zx���I�7��dR��r��h�����e�J?-g��o}Կ�S����FY�*�Dy@{B>1���s�{1�{���e�h֪wÏֱ���f_�	��s����L'�3��^M�a$n��j1Q�d,����|�k2u�i�kq���ut�ŸK�C����eڔ��F���@��+�9��|���l���RŸ�d`W�j����S:=^���X����)z�$��}��Aԫ*)�hn�+~����3�pr�/4�����6c����90����ɮW��
	�t� 8�0��JA�]���ech�G��p�ɤBm}�G)j�
�6����؅MV�CN�-SF}i����6�?T�IH��j.M�a(�NpSD��#��v�vΖ7��/:K�����P=q����y����.���n�l���!�����ۮz��� Sb��������xV[㭙&QK��Ť�՘[�K����G��H��X|"�G�!��X����Y@�����8ɣ"�!'�Un�Ü�I��+-��͉--�d�ư:��C72�M(������K�Iv�H��}Hx�A9>{-G�P񶟑�'��������/P����~e,~h��n@�Bms#��)���쯆���W��Ѹ:eP�E6H��C��Ҫ���6���m�	�ۉoo!x�6��Mj�H�l���ޅ"��	w���y�{[��U͵��X^3��O���/�]B�����r�4VK}2�jΊ���y"a/lZK�wÕ�A�DG���A��WH��b�0R��F���>d.~l骖.�4UI��R�� <�/��,S^L?<��ݱHA��.�
����.�����*�f/�W���/��#�|a����&t%	��y�q��3Z��6��,�=5{y*�'�KϦ45��}]�,1��~�9��#�=�G(N�����RyY�Ȣ�ޗ~�v� 翹���DVv,G,�&�{��!t���R����x�q܊v�t�MX���!�LI��"��C�)��LC��4TO#C�o~̟��
Y�ۘq��N�.���$K��S�N�38�nI���H������"�*�����vZt2�,�TH_-oBbh?,y`�Us���v �_�v%��{Q�������u$G8CP��8X�'��5+��x�{�s�"��0�T�"�:�ɢpʆ�%?/���*uE�M*�Vu߈ڲQ�Ͽ�!����0�&gRDa}������KS0H��]T��٢����1�p抓k��f)7�XC�u)�zdݖDc%�1���4�[����S|��.�~�V�� q4b���,9�֑����'(} !�*���� �Sl����`l�B�q`$E�'�G�d��iv���F�W��]�7���~Ў?��z��Z)�D$&zc`�,�����ˎgD^��O����H�m'a)`�|w�$���bqq jL��#&@�=���SU{zvLLҥ#��_���6 &�ܠ���4��x�q=�#�I�m��m��������$mL�����_d��w-H	����0�%�g=���s��1_�����PR&��5��W�+^�l��>Z���8�N�"�lmu�Ag3�0�y�S�|@�ح�8�XA�:�������
�����2��R;}N��Գv���V��u(�x��JFo-6�̃.X�Ki+d�,>Bu�|cw�٦x���Y�|��$�T�����E�ْ��W��#�����ܨ��� ��(�.�>��}��4%lsQ��2�z'�P�5 }$Q�� ��Fsy�!���v�����V<�\��Cn1�2;;s;P����R��xj|e~�r����L�WV-^�O`T�\�����B�=n�x��4( �d;���p�����XM%P�,[c�4��"��Ţ��i4"�&���e�a5p��d�/^f��c7Z��n�\/>Ze�T\|.#��h��uh���N����z"�.K�JX�:&~�I�U�,�����-b�4�Q�a��4h��,Y��<�q��H��|;�;���%�6����O�o�����P2�����t��]΀7>���n�bt���'�$���E���n����PY'����Tʱ��}�H�b�3ț!��FhUCGq�d�����z�s1�ŬdcvA�A)v��&��×�-�s���_��)��N}zD����S~;Ɛ�p�)�zLQ�����b�|����������A^�f�O��_�}�Ab�{:>﷮O�	��7�=G}�H���?�(q�Zd�`u�F���^]x�E@Ï` �ꎂM@?��x31OGY������7��'Ͷ��c���X��J�}���US��ݖ����X�g����ϓ� _����k�\KR�Ѫ�r�Ey��Q�����nր�	�8�m_�o�!O��$�#*:��CZ=j�1�Q�+d;��d3���#���Vd��2G�֒s;��ؼ�hG�H�~ �~:;���3����" 1&
sI�`Z�Ǭ#��� �
k�ٻз���H�z��x�K�$<��9�*��pp�q5���5��h�L���'��M/w�6�L����,VV5���I�c
��R��M鰝��#r�X�ߠ��)I�v��/:~�i"5M��: ]0��^Ԫ��RT�.Ĉ�:�gvR��d�j��׊���'b�{��(������_�,�ϧ#�[bR��0�����ѥ�U��l�R������<�q9Wlj��~�z��*ۤ��!�,% �����Jg$@6�h�_V㺜�n�z0�ʀ�0�ܥ��+����gE�� ?Q��A�!3��
��x�HHEM���0D��v^��Q^[!�2�z�߲��s��u�x61���n��q�?#rtu�\�����%�j�,����YJ�*�"�ܨ�l����d3�-�c��T�X� ��λ���qN��x�4��r|�d����hGK�2ikCD,b�p�}T����$O�*Z������
O�Bz$��k�5#[���<D��c(V� tn�S��{���[�.�H�T�tؒ%R��lO�_瓵��}i�|�j\Ú�MB��ʍDK2F�Uwl��i��j�>J43ٝ��T.�7�U�1�o��0t�C��.i�y:f/$�v�-=D�Vk�����b������3$F@i�9�@�ĭ�8����
:�v-�w4N�t��b�8/ś�M,�5%�P��Fs$��M&����!9x�=	�+Aq�ͅ�\o��b��t<�G��u&�"x���	Y����&F|�����Ok�\s!��-_{������0���=���!�E���Ҟ��M��0���$R/D���u�9�qQؙ��̛���Y�`
︷Q����flj��v� .���� ƲP�\ٴ~!�]sٰץ"k�eߨ�\f�Zj�R�LQ��D��i��y�`(oߊj9�2�������U�Qu����K��(���X>��`�T¥}`[���°n�+
@���m�!�s�t�U^��ӑt�Fۻ,��o�����o}�B�.#1A���ƴS}� �c��P��C�
8�< �n�㋪�hY�,hx��C����Z�'Pw���u�C��;W���a�b��:>B�,���tɨe�uI>v�1�$/}Ć=���mDC;�,��1��!9�s�ܝşSN!'�ar�t�ѽo�8z)�i�֩�f�\.l��
/8:k����6�z��<�_�%��Ɯ���H��� ����[,��Y~~B�Wo�tG�|t�̣PÀ��~��IV'g����U�V?B���i� 
��B� ۩�.����������@�L���n0Ϋ�l�7'��G2}����#�f���Gv�LSBG��Y����O<��v̽���u�E���]�g����.Y���]]xw��s�e2��l��b��/�� )��Ch�D�f���=z��S��D���@���(�P�����<�_��h��w��~?�`�scw	߆>�S�`P����&f �$��"����r��v�fr'���c%I/�����������/�4�Èҿ_�6�����ͶJT*�Cb�]k���.�#�)�7[[����U-�>�Z��%��L�f磺���d�Tv���1!�W�#S�T;.k��a�
w��N��F�N�4~K1��9��ח��:�����lj��=�ҫ�
.[�TD��%@*aU�,R �x�Ҧ�Ɓ�:����S��1$�q���k����m���um���kV�kO:L�C��*����.+vK�J�|]�I�������?�T��K�(�Q�s�%*��쌘�%6t��=N��r���v0�F��'P�N�<K��y,���>�\������胺�a� �H��
�]�Z���.��:nl�7�w� d�^FJ��i$4�6�b�I��zYN�ګ�8�O)s�A�9��N�i0��ћҋG�b���ln��&6��B�&g�r*+j{� �nh*q".�$����;q�iMޮt�ˌQ~,�b�EA�0?�0��t��R_��� ?;��c��ԤԦ�ǣ-�d�"W�3�m4�7"��CPgD&�:#wK�1%�ו��$H��ӡ�����F�]��g�,§q}�˹�M�BA�*P�ʀT��I�V[����4�n��h�%VU�y���6���r��n������<�FV[��'�B*=o���L9ω�M?C��A��'�ԣ@����U��S_�}r�F�_	�s��"�ȡ�eX���~2�����RY�[|*M�`�I~yJpO�V��YE}ܚ�9�hpw���և<� ^g���)�h/�G3zv�����m��Aj�ɶ��kZ�31NY�[�`8�Y_���!�6��B��g��/^�/��H�/dn���G�T;,�ʮ���1���h7��"�J���.�����H�n����r(b����pE���n�� 5���`��AYÓ.Ƴ.�ь��8�%�Ϟd��c~1i�&�v:곋k7ˢ��!���V2�|y!��i*��\}���y�1ˤ�~�#�!ec�v�s�OT�<��g̬���ؠ��Ed� �EO��}0s����a�_���C�)x���B-o��	L!k��/U�C�*�����ޘP�=���'Dl�v!����7����A1	k�v\|DTĹp��fUk��T� ��T�T
�Q����-�)!Έ��;��t׭",�x�O��P4 ����W6H+�K��YC}�0�4f�����]s����K2�ȤZ�J�:�z�Q�A�R��T4��X٤�7�lP	�	��bK�����k5�Ƅ�~ �U2 R���	a_e�s}�
a�&�N�ŉ���f��k69�{7���ѹ��z��t؁�kd@�s^f��?ھA�~T���ld��V xq���?��{�D�a�8����"��,*V2��sO�1���SdR$�%�,�h��k��p�q�"�z��d��"-U@���_'i�5H�k��k�
}9��9��H ��x�������\��R�+	��oB�����Id̶���?��-���Ǹ��|�����	�����v�i�T�#�\
�h_��Wۛ4V����<Q�ku�]�9����g��g_#{/X^<��D��9���1c𙙓���ʭ�6w�7D%������A*���1e��JQ�׌y�4\;^��c���a���c��D�{��]>�
j�'��$1�3�� Y��q��!
����YdirPTnèuCi�p	�2d���ਗ?f�4H��<lJ�������ݼ-���u��4�O�:�J�j�v۪
�'���Ke�;+��U!_�>��?�9��rc`N���ɠ�, y/�4٘t��W��_��U(P�&�ͻ���آ��
S����T�['��C��3�7}Si��_)�i���.���U�)���5Q�½��uY��K�¡�i�vL��-A�(/�gL�+���A	��R/���ܦfv-�3��Z�ގ�n �c��<.����yp�`���QKKZU�O��]P�`�7�caB�5�Kf��*��}.$7!	F5B+2����.�)�tRd�ö�,���M�-ٞR�xn�A����c�j»l�ݽ`c #x��'F��B�W�J^g%�-U>������,���"R==�h�hNd�Y�|m�у��qP[^�A�.���rh�9�Vh�g�I�N[CMH���/��7���f���t�BB�����kw3Le'�}�;�a"iM���Z@�q��U)J�by
�z�2!�������� ʘ���f�T<�pE{�=p����O�o3�!xf��
��������Y���۽_�7�d���X!�$��`=Ra�<�^-}��^�� X�_�B<8w%/�D��.P] �!7�y�J�����yBBY�ź(	?�ùfW��&�$��(�I�%�Aс�(u��A��!#$`���Y�ƈ��>�K^�Z��¤�F���8����^O@���h�����zڲ}ީ})G%;�Eh��ϲ��ժ���Gb:?F�ZKb�K����B�P��m�)8�;�U*5)G�ŸϞ���~���;IÒ�r+E��6���bt(:�bj��8=���ܝ�H��
�i�#�.�����c�����B�x"R��J�=I�n4����(น��ᷝ�kit�>[R���ڶ��~I(<1��_�-�?��� �J��"{1����(_`�4���;9R�6���Ov��Z���m�D���z���P��e]�A� �1iu�o~�7��_ Z��h|="�Á�	t�'�h¤��%l��n1��N|��L�q��S@M�����J���9���~�M#*���Ra�r�0ڢn#�pg�|�F��ĳ�`
ǫ(%�se%3�~�_��f4xs��ǎ~�YXņ���Ҁg7���Sn��p���8`D��sR������{������y
U�B<{t��|��(H:s��G��#	w�����.�O�p�Ol�����u���\V8�X[h���`���e�{����2,\�/��$L�P���tş�����v*��Df�~������~��ų<��N���T���5�2�㒌�j��dj�����@)'�S!W�b���un��px� �H�-i�;�*ʘy�ԇN�KC
�Vv;E�1�_�����]�������.x=#�39�$�3��<=�A���vt��?�)�)�������P.��6ț|�瞅�L��=�Q�63u9��c\����=�a���+�p�p�9�[G�ٖ�'Vt\X|���{	�tz��2Oʪ���wx�҅�Z�� �o�;��轣��?�O�e%��g�K�)��^U7��dAx�2:޿-�l9��=�:�������L��M�Q�Q�+��9�J�ch��1B|���Es�]��zƢª=T�X�d��
�M�YQ��\`����n��V��7�:����5�Ҋ�!���2U�{���N�А,����R4��Ԃ��� C(܃�6C��K���/A��%��-ƫI���M]v@GZ����u�QjK��})���� $��?���}���b	����ڣ�oG��M���Ze�e����[�{ԃN�*���t��E�EL���pB��Ĝ���)�*"� �G�}����pm��g�����(�v� .A���v&W�^Y����l��(��fA[m۬؛�k�O��7|�dv�\_e�p0�<Ձ�%t��A(��h��o��,�z�P���k���0��~�v��s�#(����x���s�Y� �]�Y��D�JIn^��(�fڻ�v�G$`?�R�D�s"���[�c�ܳҲ���bT�I��%ճ�7�A�4��
�=Ɲ�iq�e���8B%K�[ܞ ݼ��&\B$/\Y��*1L¿<��y�`֟=pGL	ѪzB�}o�R��8)鿞��D��BHɏ2$�Y���N�O�S
=޼!�^���:������ �� ��S��XoyYA�T��a���ؖ�0p�}p�R�j�$�QX\�u~*����T�'�Uq5��'�q����w{��G,�G#0�^�	�@箛�&R*��į쮂 �� u�j��&r �Y��*� ����ࢹ;i�T�_"6kʒ�$�z엁"��hcj����9�+�	�ä���?�6�[�"]�.r�V̱n�6�U��p���Ѿឥ�5�uBv�5)Y2������ W*~+��(�]��Ss�k7����z�g.����
qZ�'��c70KO����л�""�$d-J�i����KZ `g=��&���T���p���S�?3��&4����ek�?9��c�c沫�������[g�l��y�D�����sT��B�y�Nk	u�⠃�	G�V��EYT�r���"@+�u8�SPc��}w�Y��*[�o��>������/zP�b���ǿ]VbK�Ys�/$���U,���I����7��yt�bÉ(�4T�����;����Y/~Em�a�_<����\��>6�	�R�Zu0#�����5��c���a"K��{�������4���d$Y�pF�bǭ4Ia�F#��b/�M�?�@=��Y��C�g��8���؊�E2�r���,,�dyR�������`J���[<���C?��rsd����8k=7un�c��f���::t�+�4�.J�sn au�	������}��L��5s������J��B���yҐ��%�}�n�fu�W��z�q69&m)�7"��Z��	Q:	���UB	v�QS�H	��9���,�LZ�e�Eڊ�X�EV��!�?�@ML�>_e��L���N��j�<��$��`a�HT�S1�za�~񴤭�[��~ rʣ�#ׁ�ћ��׫�c1�L�x[��"n̓	�p;집G��w��2�� �g�������dLס���(Vl���_ƪ+�.e�q\�V�p����(��WGU#y]r#د�9����9�f�&p�����7�C
��C���LBd%�aW(͒���X�T)L��ի��K�J)�*	@=��@O�G�
F]�@�7���s�2�!!?��J+�\m�?3T_-N�͆���S�Nא����e�����{̷�x�J��@����V�8;g���B�lyL���%-�ƪ�t|h���
������x౏��.�A��wú���q�8m������Z��u3K#�
5��: B�n_W�}Ǭ�T���Q��s033�������-[��v"gQn���8���,>K�_':�n�d%P�}#l|1U��2��bԮ澷���.�Im����́�'�<qY��ѥ����s��e�ȜXR������o��,��uZ�/���i�q�������BMT����Ƞ^Q�^Fi8��"7���?d~�2p୦ lfD�]+W�}7���6�	� �}E�Q|����٩� ��;�t>	-~�&6+��('g���˞6C������!H�
�	yl�X̧(le4�v��(�?��C]�A�=x�+P?��<W�"G`���b��6=��A"�бZ0@���zE�dZߞ�Ơ3�\�� ���4��(i�|����hw��1E�ŮpN��i�mn��j��@4j�Հ6��sG���4}�N�������|"�2���w3&��Ҩh�*c~�W"�8�z��r��M���c^s_���4V�*U�f��v�4�x��q��%v�Mej^߈L���<�(��,ؘl�(�k	�*CM�aT��Y��!��>�N���}3z�Q�>I�݂8ϊ���S��n�ė
'5�͛R�o�t�ݗ��tQ�|b�������E;q6$�t�X7�c����]f��Ho�Z��1S�ZT���ϝ�Iy�>m��$��yU%�vG�+ �e���/ ��<ʍE$��u�����J�R���{|�������8��~{l6O��r&�n�t�_��F|_=�[f#��!��2��k,�2��c�:�b�Z�1>��?@������VZ{�t�Ã,	�z����=\�Ҧ�{椇��D1���s�W�_����㭠���`��2R'?.����̬�	0ʉU�����}�C�E��"��г��:�;\�je�Q=�?l7��(,8��ܳ����{ku�Y^ya���K������S�9�"X�,��)��_]
:���]A�ꑒ�k	��nw"LA�f���<4E&.u��C�`�#�o=Nm�U��Ȧ0�05��b�m
��A#������wo.�>��޿�J��ؿ�#(B����.��C�BgsQ}u���|Oiծ-���}�wM@lBXy}�,�T���yB��R~7�")M���a+]���!<��p&�}S(N��B0� �;9W�}��k�xQ��$@e� ���`o��*{F�#J>��H���_,57��kT�*.� ���	0Ʌ�z�9�w�w{.W�2�BH]QZ�x*�o�ǐ�r'ì;J���S��2��(�$��su�Uxvs_t�lM��d���y��RYB~��Z<�;�mn��璈�6i6m��σ HX83�ט$o���_7��w'�x7�t�!e�F��>�]������|�CB�_G��w��9�3��&g+���VV�~�={��ߞ:2�)	�ߝ�7b���2NO����\@c�#���tJo`�%��	`�#�r~�`b[� �6W�ƘL�X��v�Z�a_As9���yz�i�m�j�9$kݔ����M80Z� N����;>��"�����6l�jڸ�S����Aϲu��H�����z�}���r�1亿�ݧ�#SM��.ʲ�V+��g|^��r5���c�[0���ߩ�y0MYǮ�;jB#9��Z�o[�K��R���@:oAp�ڰ)y���r�4�$ )u�����ӧO���GM#eV��m��SCX�]�����T�f�F�K��'��am�M�F��X�jؖA���L�m�<Lk!7�ک��`&�kH�,�K� �$]����{�E��B2�n��+�5�7m�:�^ף�[�H�iƊ�q*��uV*K-�M$
1Nu�{QͿ��P�/$��!1�px'����D4�}��X;�Ɲ�F��A�����v\���qg����1i�Ύ�-�Q��p�~���smp�Я�C�A�����n�aU�����3+h�A߾�.�6ߑ�b��hi��f�{C����R�{rS����-m�ӛ�w��s]�=�i�]޼�.L�^��2�1��_bңi����D|91�8=����Te��GmR$�t�6��@:�F���]U�#��ZF�-NR�nTt��s�4�.`���]p�ab}d��?D����.˰�E)gT��p$u4�l���oG!{�п�q��[�}�&XĔ�zR9%P�xP�����Qy�S�zW������Ch#(%eM	�*<��W��q��\�z�j��3��td�gYE����z������}1K+�������EKǘ.���HT#U ��<ط�w"�������M<�O|�z���H|�yi3ñ<a����')J�im��Z`d)��V�R�ŉ�l[Y�������Ⴒ�)PĽ��dѵ�+R�� z�Y����f��z����gUCI} �4ߋ��]pǜſ��CRB��{d��k�A�	���hJ���(��JH̼�+=��<2�K�$o�	�u��g�V=#Ky�J�Q�y}��N��`>�A~���R�^F���u��O��ud �C|��i=u�d�p�τi�x�'�w�Xm�����a4R9��Wv�d�$ã��+W�a-�l�����w�h��^�Ԇ�Ѻ�����7��x�Kp&Ȓq��w�{�sve&�4���=lr5�'ߘ�O��A������b.��L���,!WD��)�D'B]7�r���Dv��x���.�N�o�4i��t<D`�ݱ�h�(�@�7�����Ul{���:�T2M;[��4OI��k_g�C�����A$�E.Ĩ�
���&��Y=���렎[~��y� HK�sg��9�FTq���*^�T�m��@�������Zb���B�Ƣ��/N��;��9b5a�08N��>�y�)�%os�ωҐre�d	�FXy�����?�.�{��IA��Ù���� _������>�FX���vG�6��M*, �,گ���][?np燎�$D	�4�T0�j�Y#�be�ŀ��N����`��^��"�}?`fU2f����R;��6,!�}K>��R�ly��bxAL@4~͍�,d�z����ٷI���|���I1-����mbV��sV�v�J�\�۟�ԉشZ@�$0h��W�c�t��m846>���=z�/MS�%���yĆ�Kq��_�6�6�ZK&���Ow�hR���&z����#w�O%t��q��(����6�>����9oǺ4h{��հ�Q7�u	���=��Xκ�ų�T޲�2�?��o&�?ڼ�S�q��\�\�U� �%:Q�"m*F$��t"������ra�t|����2��t�Y�с�(�*^�G8$isݐ�0���D*e�
~o _r�0[�NZ/�p/�pr��3sB�8fM�b�]oL�@���"9`�bjj����W��. ����lt�/�c��_�d���ϒ(���+m'5�/v��U��-V��*��Z-�~pbK� ��;�%��Z��C�_���zfV��}L���U��E��*�г*�����4���+���ĶA�.&0X��D�n�U!�����k����e��@UK�rZ�w��U#<��
�8��U^��6�!~�pOL��𩑞WUD&j�J�$n������ܽ+�Ӡ M'5�Xܜ�!���*1�$�� �U<Ƅ�D0(��Q�c�\��`�������"�X~�y��*�jd�r�1�|�n��7�ӌ+���������(è�Yܴ�܂���@w�tʱ�xݷ�U��v/����:T��+`�M����]n<|���o�b���%JI1��x��׳x�Qa�'��+���&pʣ��7�
t�4��]LC5���l��V
�E��A�m�-�J�q��H�ZL��������=���x�V����E�_�M�:��#d�w��m0-д�G��2h:[���Ϣ�~����1��&�� �x|����5&�����>`����:�6��>��7S�ޣw������`T��8����u��{{��V�;ʔh��!ӷ��2Z� Iᘦ���̥r�~SJ� ���,�'�R�G��(�{6b10
�W��!��������
_�x�9Q&(�FV����U'y������Ӳ� g����W�����؄�ę�*����l�e�����cb�.=`��uȅ�%�$E�������pgIJ�~�\�7`�f�ZO`�h��5'��4Ξ�B�A�&���Th�����[�	�!(c�V
��l�������p�s�s���������~�I�l-�\��4�V�6&�,��(��N�_�p�C�i��--����Ȕ� A����\����;%Z�B��xq�,3c��A�^�0���}����H"���d��<<�"Դ�Rg('_g�"��r��gN5����g+y 4��hxg�J�Q��N��f�4.ER�4�Hg����4%�G��(P��@������3��R�������b�x�I��@��Y�1[���O��E["�Qn:U��r, ��:F"��"�wD&�W�?}?�s�;�~�����4J�X
�4DS��o��F��K$������3'�9���w~�Ûtn��,�'Y<�\�m4H�n)1VMk���n���y�g�q3�1��8��`/��d=ך��
�z!�6�#�����N�"�a�*'�����%Rh��J�k B�!x���|tv��(rT;Y��Zk���Z�̖^�櫿��x��\�7�v7���$�kf�FJU��#*�6���l��R0*w�F�-n�U�����h(^�ik�x=�d<�`���A�,51��q�Y�cl�J��Ԥ�#w��).��O�����T�6sv�$��E�:B/^px���<�d��9�Pq�P���?�R�������]j~����B҂73���ZSK)�U�X�[�����(9���@֎�� ������@w۟�]�̹�k��_�[�%�UO�Y@B
����U$,�!~�d�S�Ej��B�b{Fh��v��
<�Ѝ����W�Y���>�&��Ԓ�\�(�����$�YR�Fr����R.Y��HUn�m2�Pw�3���W�=._7�6����onl,<���5���I	K���$%���Vʹ�4�$�u�Y��$)��"E�utPl^i�vN��-���w��Y���9u���
k���xZ(b|�� �����p���w��{t:�e�X�\��#[s9�����j�P���^E��9��g�|�+\1�u�lt �ȡ�O��:z�(��V�ȗ�y�9(E�p��qɍP�����ţ��禃X|�	^2F�VV�5�l��H�gS�nv�-�6���N >�s?|e;�o�KV������6�m�g�2�`p�{iQ	Z&z1XIG��p��:%EP���I��B (�����������,4���NV��:`x�XƭOu�晾!;����3U��ɀ �+Y(J��
��u���e�ވ��^�%�ټ:|�̾Ȗ��"�?�k�������PL}�,KJ�;�븕�;,�2���O�aS��.-������
z��W|����֩�e��d@����<��t?鮊(�kը�!=Z&pT[�0�Q���sX�����I`��J��@4�H��Գ)�#�ے�r�ˑ�P�ٽ��1_���yG"�J��o�r�H�-5+(_l�d#���F�>�Ӿ�9�>9��ܮ���;.np-n�Hm~I�� _��m���R���!�e�����,KH��1=��K����|�	��y�#3	��s8�7%���������}x�*3;$ �e�ۨ`�D���[CV��E䄦�U�1]��!9���69+Gv.!�Hv ��Et�'䬄	�]���>w���-_ �9��.��v����Bö�˚�:{�uFt���
������2K�o�yi���хB9M9�fH+6q�)�>�:ɏ�y%vU#�|���Õ�İ��I�K��+P��qء#L�z��밻����W�H�*k)7�����'�p��Ca��,�o{�� w�x'<%̎/�|v6�/YB򜁥��r�o�=���w�Y�`�)�-5껎2b�J�`̖a�}��ȴ�|V;��XB�[_�̍�&�Wg��pFo**°�|�ޝ�oBr��niD��l)�9�ŴL�Y�̆U�s�c6��*	]��~2��S~�|_��R�p�=��J������`��2����~��B���]�=P���z���8�y�r���nk�ђ���K�� ϛ���䤋�
��AB���4o�C��(�{&�2�08�߀����P�z<�7���C^S?�a]�[dcc�ŀ>���S^NQe��~qkn6J� Y�����~�O���⹗b�=�����wZ��'�W�o�57�>����<�\jO� �;z�u�����F��9+&�ʥ,q�w����MkL����)�F�tf�6�Ʋ�_@G�[��({6d%��o�{�����la;A��E}��2f��[fh�����}�}R;���^K�\Y����ۓP�����Q����8/ܫȆ��zG\�<��M��[�uѤ�f㱛o�D?��z��>�n������YS 9P>��:n��	|�0Qm$[l��.�u������� �:M�@�`̻���+$���y�C����D=6�Rػ,2�w1�מ�;�N|58wq�S-��o�X��TaK�7�jk�;.��@[/�f"P��a:!�򣬫�5�)	>�Ҷ�E�̯Է�"L��!�v{��1!�W�#:���(�B㭞7BR�}��ة��ݶ�dV����b���
�^�h�����ͽ�})�ͬ[��㟧�x�Mj?X�ZGq�dQK�Gݱj,DHī�: p��`�O��d��cՔg����,N�}]�$H���5�/���4KI	�xi���q6J�{��4��a�oFb�]��^��w\OU勭%��	�NpN�-��:$��yU�8J2�̔�ѩ����5��uT�H�F��3��2�/C�����^�Hzns��`Rr%�Ig�q0��:�Y�w���I�.�nĿJ+oQ�P>o��̝3{j�������)�/��~L�MPa�2�����"�,�ڭx-t������˿X��7r@Y��k�ǎ9Й me���-E2/Ɵ,���& ,<��~Y#�8��-W� <�8[��7����R��B�@]&���-��Eg�G?m�(���}�ǰ�<d��6U�f�S;����"��I�ԥP-��o�Vv#+A��͉Z�/��n�mh�#Xw�bXX��N-���Cc�� �p$����">�k��]&�-@��#�����Xc����6"s;މ�hH���@�����t"[��IDւy\&�T[��i���ˬ�I��@�������w��9��{x������6�b,��t��mr�I��e�/}�Yfs:�� �ޱ�QYe��<��D)R4c����ádH�d��Β��գk3g��mlt=��o���3�OSc�Uā�c���$����Ņˆ5��(
2oXb�4�-�p�P<�J�U����Ő{i���i�R��y�u��9�(�r���d͚g�n�!Rڵ�n�iz��K�ң ����D�}OÉ��Ή�Q٠O��� �v1y��,��j���a2��,-��ȥ�-2�H�R�v�(g>�x��F���vv�����$S��f���k���	d/z4�����쿀LW:���,L
��J�d��bW�Ş���t>�e�(�?��v� �W��}([�r&F0��q��A�M�1c6 �s�l�f!��\RF>�x\H���B��!�����,|�W�Z	]��/B[sM�~ ��̒�����|��a����z���~�%h�|<��A,�H,1SB�6�[}Fi�^���	�X���)H��x�_}u_�@������, йˤ�l6�3	ħ�� #���^ B��ȁ�����*�v��e��F��r�&�"�%.H��5�p������I��K���ܾopӉ���/j'C�R�(����<�Sf�,W�']5&ٜ���0`�V���u�����P!����Y[i�ۄ��+@':�hJ�b�����D�N��L���e�k��1}�\E�6������Ub$D7L��L�`]�T��^'��g�p��,����#��R�'uv�&�|����^b�n�P:q����WZ�$邉4⻉�ywz�#�OZce��Fz&?Ҭ�R]��"�K�(���q婿��\�A�$~p%8��W��%��*��� �a�좬�1|IO��:��������;*���jssi�	���u��-�gtΔ���F�!�Jpx u�@*ˊ��+����R���ڀ[c8֔�v!�`\v�����}�7�)�q�,������ᯠ�y�ZZ�=��+viD��B�)�x��m7�a� ��@�H4�eÌ�*f�i�j���ؾ�r�y�7row��/�T���O�_���1�y�	�����f𹢽�Gڝ3-PIhNl�]��#�_m�tW����|b������C ?
����m���VF4�%xE�[�~�<�o����ǋ	K�↙$w�3�H�ӻ��pRHݗY���cZ[�3��|��uI�H�]�N��=HP4�6>�0�����>�<�l�@q��FJ`��*ٓ\,�WhrFf,�:"�]�A,8{�=��-.�1�2��[�?w�$�od*�K���	.�u�(��D��!(��w&������;���)�3;A݊{h�/���ڇ����V�`�T�~��LO#@a�^��ϮR��6��_Ӊ(���e�k��_^@"r���?8K�h����X5��Z� 	�ApZ�[F*��5���FM.�ҡ|Ο�N}`��Fj��-���Jw)��KagB��O<)��kpT$H2��#�@P[`�9sp%�(��o���&�j�?聲�_#�$���z=�T)5���#%��2w1���H!��(o�t<1����{85v5���<f@Q��m0R�m5L[�5���x�#̅i��$$�����g�,���U,E�{֨ǾJ�?J�7�0ZR����zWSV^�o����Eז�'%�_�Z~�Y�׽Ht�
����(��P~�������?��5�f���� �nw�Y>z��,R�L����8�ӡ+'v
�B��Q��S��C�	AG�W��C.4,�~󌦳�$�=�p"0j8I�J�2�1����:�iW7�uy�qB�p��x�@<&sM�Ǫ&7"o���d�����3����X�!���E#B��RK�P��L�'���I�U�,z�#�&n�K���[дc��v'��8��O������j>��!�586��Xl]0Jo"?�*����:\�Gs�C���pe�w�$,4���]r6L�C��g�� Μ�N�%�Ҙ�B�(�*�kJ�}�k.�-.��z�H��hz�J���$o~���d������n�K�~v���:;bj#ݞ*QnM�ō$<��Y�ϯI�!`�쪥�#w�ܒG$�o0�U�,��up�Hx�Zz�89caqUBV�ݬV�rE=�RNy"15M��qQD���3���]t�L��9��!;���ufY��a.�(	t�����s�L��zzUv���}[�d*����������b��ik�V��g���.1�p��R���ś�g|5: B�\���	�~�t���!x1�ٳ��S�tQ��?�Z~�?u���~����X,�R��g;&v|A������"��Q bk<R��tM�Q�0���K��W�9��-BZk��>��MCr��a�U��o���'}UFF�ֶ�r\����D�:&���%R��9#�zv��ZNN ���[J��&�xf�&�Ne��o�Z���HW=v�_f:1���<�f���H��|����?�#;�F��C1���/�LS�,���&*����\��*��߈xoP�����#G�'����ċ��B���2�cZ0��3��+�KH����\5 �����r�)VpH���b�Re���6�sIlI~2��$���p�=%�aի����v��C����(�+}XxP���̿K���6�1΅�����>*��<��C�Uf�jP<T�ԁjeԼ�t��k����aq����� �AY�;k)TzK�);��\6�BO�t̑^���[��?o`�J�@v�B�ՈL��M?�=d^�� ti�v�`��,��J�I�;�G��e*��u?��D�i7��f�BۊIb��{r��	ft_W��r�=�-Zt k�"G�"��R�LSy�ZmϴCy�?�������*(�#�����M�Ɉ��'���������/@�7��j��Q���򸙖���n��rD48�ā�m{d�{�bpǋ�����O��]��k�uH?������Q7��Ԫe7�slu���tJ�l>��x�\1{́qj,�.����!��
@���^фX�U���Ž-���%���.��9�)u�?���m�J�>�\���?��l�8��&GR����S������9�xs�����ç!�a���'}/�ނ��rӝ������T����&�j�W���q��6�X����%ר���+�麴E%K���@�iv~i�u�0���/����%��W�HxorO�.J*��H�l��:Wt!Nu-j�씸�Ï�0��� J�6�?}	��0J��ki.��ѳ�+]k^ٟ�d��T����=�iW��Γߛ�u�<�?�}���.6H�hDY�NL�=�l�Y�McnSyu��Q61 %k$u��V�x"jM&w�����	�{BX�<B�Q��ٴ�2�ya����屫o�3E]��G�:��.aIʭB3;/����:I�;�*�I�0�״��ŀ�H�cjK�����Cnw+�/�0�ArA$n���O����>"�V��A�ߦA�A=ExeX3ݭ�2�T�>�ë7!�<ه�ӛN�O{�:-ѕ��NT�쯥t� ��un���{��#I���ˢ�5��8*)wVq_��P����t��ƿ��U��|�6���ƺf�:./ ����RP����W�q�$�Z�喨4O��u'���k'z�����S�מ�y@�Ol$�܉�6�w�&�k�Q��ed������3N9.B���H����%XJQ�g�ǐH���r��X�m�$"Ou��E��i�ܸe/A�au���J~���Q���>k��T��mtNr�D%��4t�[E�Q�B����!:�M�B[-��U.���9�����u�u��2����"�v�{d��sy��}\���%n;O�]�s�":*�]�#���N8�!�g~�0S�94���� �T#g���OVb%�y�@=��.�P����Ө����Fi�B|:٩�7���C3�۾"��c	�nB���������_n�L�pS��;����U����sg�:�eJ��|DD��O��������S�|��X��>�5�!��� Gq8ҵ0Y��3D��j�[�T#�0~;�~��U�"�F6O{c7��2X�t�[�Z��[�畸�<Cb����l^��Z�IL�g��[�1^�7��%@A���
��L�6��c��g�I�.��%J���,mV�&� _Ѩ$b�n�X��Y�@�&4y���/�֘G��4�đt���ý1���A<��=0���9}�	Vr/z�a�CŎ�ӹ�@9Q���o���(����5u�=
��l$�7���!e*`L�a�Hg̪�ߓH�r�I7��*������I�b��������>#0?ʸ�{�=�7��:P͙P�E�5�ڵ�=0jt>�?Ä����6~��"�K�>����.	���Y���X�/4��מ���n>ōU�7�t�B�r��������c��lJl�-A�-Et�58�v�A
| �aƕ�����8���р��L@�I$l0z�t���<s��Tq0)F;�+�:�r!�?��K-nxԩF���d,n�]mf�}����]Bh�r�Y��?�{(���Z?�E�c���UۊI�i�^NK�oM +yB��4Lv$�L����+�<�\w��V)�r`b1�I%b��V��ml	[����wlؒ Y.��X��lI�@�,���	!��>����9�
���0o�M�k҃]x˧������P������Ռeb?���~��(���ݪ�nX�t8�f��(���&X~���;I[�	�N[KA|�C0ڪ��#�c�sV���{i���a��yA�_  �GsYI� �\�t�c�(�`9�8_�&���C��yM>�6��
�|To)B]�]�Ġ���	=����#=3�G�0���h�a@M�6���K��fC�<��B�;�C��ٌ���$Ls9{�嫧͡�Z�t�Ē\7K�(�Q�GiL@�3�z�8��I�3h�ف�"�%B1�@*�璪�2jQ�J
]TT��ޕ� Pm/�7�]m�K�h?.���J[���>O��{@T��v=*{��GkrH�ށu&��a�5���0���Q�_HNu"D���P�n0ΰc���CC8��(�֨l�b���-�
)��Q~��5�D<�޶˸]&�2
h�����ix~�$2��(�:'�s8���0��I=�W�KĪ�pSv@D8L�Ajg��'�~�<��^�7�qG��F�}��֞�nr�S�#�_��vHy�%�Tjhs��e�|�;���u�S�X��M��{�E���9߅��1��v���H�.�@xP� 
M*2vG˿~�/�m
������:��"�6�k���s��LJ&U1))e;D%���n����HY��uFj?<}�,�2MUu��}��˿�������B,kq�KE�b�ӧ4��ʙ�ze1Ԧ0��hQX/���C��Y�tv���F���~:x�� �x�k��Yǂa�hQB�i�yu�v�"q<�nx���{��W�Hk$�H]
�����T�!��1�潕N����2��2$x� ��'��T+<;kU�o|�s���SWR֋ �T/`��@���,�ϴDE�E�?q�p��a�'p���A �?��w��� ~�o�o��p�-�<H�w�{ǝ��kt��呭��^��,���∾A��N6>��Sϡ�]#�$��sL�T��8�Bs����,]�P0�i�0���ip���̄ϊ|��T ��ڐW�"�:�y(��ε\y17G2j�';�q���Y�4v��p�>�*#졡�=m>!?FE ���{�������m*��k'W��aV���w���	���d*�fD�,�O��MJQq�eG.�[�i��@�@���Nv)e	��qOtw(�{�]A�A�I�'?Ԋ�˜]L괰ࣄh�}��WX���RT'4�6(��n��f��\����
�X`#zi��߸��	,4��"O�Z+̓{2=�y�A"�dM��	2Z�X3I��s�u�:����M���/�\ϵ����v��Ѝy�"��(Ǫ�7V:���P��I��U��2-�($���,Q&kD�wo�N�6nS|B����7��%uC�I�i�4�G��򬼥����tc���/�2 T��o��q��4W�(��pUYI:&V?ڻ�"OE�
h�oU��8pF��C�?q��X�|�񅕓U
Y��9J2�.V�Ge|�CޅJ@��d�M`bWQ(����O�����3r#Ԗ?�<��a�|L�9�%>N�/y��nl?P��?�4e��{�,�:�A�l��k� ]#�\C���ﴷ��eC�Fo:ohR3��?5���p�ڵ�t��hn�/��QO��rS-����A����:@2�AL}�`4�Iզ�{P��yE!"�+�|��\�q�J�	�RP����{�W�:	��#,:�Q|
�J�Y(�~�`R��U9*��� ���#N��1�|�G�~Y
�MJX��o�u���F�($鸭�՗n\�R�l�B|���䥽��n�ǈ�q��6�It�R��أӡ��w<�+����_���X�TA�T�|�N��W$�/�^����E+@�5
aO����Nwg��$�S=��V���\n��
�-^t����Y���mɞ�!L?v�Jnl���i{�[��@�V?��B�ܻ�.��:�A��[�ULnRB�>'u�U��XY��U�_]4M���~KD�@���Ʀx,�`+Tϼ�D��!Xx�,�1Ǎu1�dUrQAp�D�%��jK9Lذ��)�B<�w����V�Uq��r�Uc�@�C9/��M���ə��N�Jr#�<3�|��1��:����\c���y ��l1���\5������!��:�����Vcf<Է��0��"�>�`�Y���v|�n������o��I�տe�{Y)q,�y�#�Z��p$��Jt����PJ�}w�oA)�aqqטi�82�}\Cjq��c~m�nһ�{a�F����M�S h��6��4Т�����r�-��{vt��_���ʜƄ�M�\�����*����7�߄ ���N��Τ=4��~0���\}�H�+���XL���ڟޢ�aS� ͫL����O
=�|��2d6ṳ	���:�N�~��H���#�Vn�묶Ԕ�eq�
�XuI�iy�N8|�d	-W���<��k����}���k�2o��,(klfk�9ƪ�=�)�R�~ʁ%,���$a[˼;�����@tعMa��F2�U���������YF��H�D��a��ބ��ZkMMgb�&k��4�/�ʢ<�0�k�)G
�� (�i&�?���@u_5�!��� Ȃ��&r1�����>i�� x�������Z	�J��z� u6�E!a��f?�`֔�Hw�B��g���l��?�Đ���ܠa[W��q�)�0IO��ޒ�`R~��Ma�eh۠���
��ˑ��R
��M�G�����8-�J��M�?��V�%=�l��G蒻D^$	�b�J͎0��m4��k�|�&�*��g1V�p@a-$@۽Ԝ	`\�,$X��3�����Ɂ7�p~�?k��8�!�
IY�[��\�zh�ӕ���4)�<�5�����Gc�`�e8��O�c8E��"n���V��n�=���nЋ
T�Q_���������>`M��92l��n���j��I�E_0>!:�dLf���C�i/XD��a-�L[���_"SDp�@���F^���?��G������u�Bor�:ƥ�_E�8*M1�6��D��.53�ݞ:��/�|Êҭ-��h�E���(�Gm�^3=��g�0צ Xq�~�b�mco^^�#Mf���VM�D�\e����S���+_���3̣jKQ�2��p�W^��{E��^^����vކ6���#�߸��z�{�Q��)f�KЩ(�|��0��l�D�!��c�]l 8�f���0�U�8�I��$�L��Lg�z��=f������k����h8����c1�ҍ��2Щ ����,-=b�����,Lo�+���0��
e+|@�&��-J���4�������e �)lm�#��0�m�����P1��Ѱ�!�NEu|0�#4̦��j}���S8x�ZďA�ˏeİҡTG֩����'��IL�<Ҩ�¦�ZV�"N0 �MxùMIz8��ۮ:��_o�<��W߹r�X�4p�G�,��8.��,yZ��{/����_Pn�8c��h��	T\��2�O�@��)ҳ7@g��Y�Ea[C��ٔ�0��k�=7��g���u�-7"�אs�FV�O*%&u}2�;n�E�4E���⼏j�ބ\�7��O�b��A�?�T*�n��X�47��g�jj�=�ң�����x4M�8ᯥQ09��%��b����B]�l#q+�����#}X'�.��Ԓ�)4�m�+֨~�|ӡ�/y�*�@�lc0Q�}{����H��II��t���{����~P�"�Ǒ�i"�{���0���	6e�t���O;N֔���beeyD��{Wu�����.�Px��&JI%~���W���%W�`�C��Py�a�@��Q�A�	��ܡ��6�����Tp�Q1��#O��IR���G���U��F���<�*�@$ݛ�����Wg_]rߕ_J�)"������-����Yԛ+��^!�R��p�|�|<oy��˩�4��P&b_m3S���O� �u��q�v&�-�EP��]��r�f�0xp)/�)~o ձmi�����xH|>��~�Q�]�;X�(�{�w:�ތ�IĈ�~DaJ���+_��4�[���"g/�D[������W�9ħ�����e�@i]m�T^4�)�G����k� e�I����F9�׭6�kg�0����.I�a)��Q�b��&������҇I��O)�f9?'�$Z��*j���j_u������6�B�� ô��a{{|���n�!�(�8�A���UM�y�����
��O8��#y_�!Rdݎ~�5�NZO����96���HQ���޽N+�Jxo�d9HO��!/#�"�\�|�g F�(4e��n�'kT9j�+��^b}�R1��e�z�b�x�A��������)!O�CRa��bsX
n�!�Oy].����d�)�!�c���_s�ߜ~���v�S��2�����]�J<t�~���h��"&KY<�P#�o�RaDVp�csM&��9��M��ߚ�����N��^��@j��D�O�2[�P���^�� ��or��݀��1Wx���	_V���.F�m�Y0��q	�(<��mFzG�l�p���~�#س�R	.Z�xB�fg^x��4��O���V$�(��OfL�;�ڗ*�K��}�
aV����F�`�����/.�#��pY��Y�j޲j8Ȱ�Ql�mD��66���W���Ɲx�o2��fL9����:������U�6��<w)�/��g���];H.�Pfb��-��kSlP�����+�.�2/x�f�7L�W~�=L\D��~K��U���ԓ+6�	>j�C|�_BV*�EMc "����^�3ΐ�b�t������A�%����Y�Ҥ���ъD�jR�϶��K뒮��ޏ�/|�i�w_/@)��*�CV��ճζj����P�`��'h�I�n���c��m���E�A��݆�Đ�0��o�^���l��8GM�()�>���k�+Ul��v�ʺ7(�oh����ɚ\�cӝ�e;���`]& �E_}��jk�� �[�S�nZI ��d�F|���@n1�}����w-��ź͜v��̰��v��5�X�o��чEQ�Ë���
'�p<���t-{\?�*V�#��Te�/�<=�PЗ���ǝ ���f1�`������J���/fs�¶,�����	#.E����ק����Z{Շ&��'���W�-*�X�_C�D�q�=����m�!8�y���_�quU���	��hE��6�Z�4N��vP�֕X�=�'q�+B�k[>�/�VlYW	�?d�r�"�~�zە�(�s�m��2�Lǩ�iN�S�c�>ǎ�g�1��2sj[�i|��(z�uh ��@%a�����,
��n��#����䭾#����Q�����	�;5F��L�ֿ�UN]�0V���f�7�-'9��bCa%$���{�nU���d`0�-O�S���,漥���zy��?�e�C�J���v 5�>d��t[^���M�(�߾hE����.����~�D���ߘ�] ����ف�#IH��Mp�S�'lsv�D08�	��ױ�M8<�3��v�2���M��h%���Q߆�VW��I��k���EF�y�t{����/�X�tJ�w��O7�Y���.@+\���쓹��]�5�+��U�)�}v9ʬ�>�������m���q��u7�-6���dϠ Q�w>=W5D����H=o��7!��o�c����;{�%mF�����r��?��;Zw���R�9��m�9V��qVV�/Y��V��Q�ji�	��H�[jВ���\Z�:c/�v��dD,�e:�R{l�o�ɔ�Pʊ�j�5^�w�d�S~�x,J���.���PM�LǞ�`�UA�b�� ��|���)rT�`�����B71�՜��bY��N��8�>�<`��p?��( ��;���έ��kjR�Oj0��1J���AVZ��?��I���
o��`I@ǘ�q��Qp�O#���:�����D�g��݇��! '��}vX�{V��u;ߥ%��b�{��9��W�.:��6�:��b��]��YN��;b�u�3Z+~瑿��/�X�bZV��گ�&��I���;�R�6����q��_r˳�����W�r���q����e+)�;�DA⁃�:|O'|]�݃�~p8 2e�Q� u�H��>���Q��$$G�錣'!�/0�%�r<�E�8�rO��(dƞՐ�@!� ��i1���u�O	��viI����"&9~,@��1jA
Q�=�&ه�Vr�f3j��T�ө��Z����$ -��Cr5��\i��a�w��>�����,3K��(�W��G7��[��Sqp[�U�]*6(&���&��;�B��B�%��Ǥ?���p}��v�61�X��a�u�א &�{����򝙊C�n�A�e q����lJ�$.�O�Ei�DK�q�4�R��H�&cJ%�
R�ʾ�JX���� ��Z%R�RNe�
��+���~���	C������%' &#�j�ځF�p����P)�3b��:���躸��!v��A^n�/1;Y��y��v@%g�?�R�V�i�B�1���B7�0�Rl��B���ab}|J��n����Z��ZΣ�xm�C���W��닏�o�X�.����`ᡚ�e���M��ވ��`��YW��]l?H��{N��
�eo�D�t�@#W���=2R�Z�>,묃���{�P�f�j��]��fo�*���Oym�n0Ӹ��8��s���^N6,рE�eK���c-,	S��r)��vCc��(�$��&���>�43�x�H?»o�E�H���<��ݦ���w^�}:�L�ln��sy��[��[F=A�cv#���AW1l�Xdؾ�!�ʻ�j�Ҥ^QU�{p@~���z�\h-Uv�X��ZԼr�����R�w0�N���"�����^��,9�/��!X1�i�DS�~���FL6p�ª��;P���B�I���u�[(W������gkaS.2`t�.�Yy�U�9c��xmپ�����ڍb<]�m�������[v!H���7X�����)�9΄�,��������Sh#��?����S�-q���{T)1*�	d,3�����G2n�Q�>�N�Wԡ���3T9q@��!�go�i�����ڒ�hz�oo������{��>�,�Z���u*nX�ID�h92�[	V� 6"h8��^�j�U��՝޷�ʒNf\�m�G�?{� ��i�@tFj���vB�#J8��ܰ�w��"����%3���Tj(U���j
��t�̦����Ȥ�cA�
���'m��B�1jk;��E�r���AӚnu&u_���߽ȗ�а��_�,r�;K��ᶴ:�&J�����@V��ԣ���r$�7Cwp�s��lm��Ɋ��e-q֝�Q�
���_�%q��%���N�%8���p�~l��&�UC�+�jn#�>�k��̓���O�̹b����ˏ2���<;�,�a��^���9�� jΰ$�n?~�3����B��H���
Zn���W�w`N |���h��q��1�a�c|��`?.}�w�Rn$.>�ҕO<�ʸ�XCE��oq.�*8��R;�r!0n#}.�_���R&�-zˈ��ֲX��S5��ي,5�8�t��o#k�#C��7�;�B�� �|�q0;����:����N�_{XV��Z�bv���G_ '�%ʊ+��u���J}1Cz�����DEdlu3 Ku�rU�[<��vv /F��]Pwdh���}��R�)M��M��4���+ї�����<TM��'�*�E{���������|:���Ӓ�^95h/����2����@�V&�����bT��GE�W@tyk��m\X�����\��x}�Ϗ�r>����+������F7�l����8��r�㠠��g?Ʀ׆�I�.�iD��b���c�����"�Z�a���kQTݧ#��l�ͱ�&�]IW�������*��bDB���D=�S;��Dp^��5e$���j;�3����֢u]4��ÿ����Or���y��i�2�N�b��'B�1�J��$��dn��8z�G�+�������y��D���h+�'¿(eB�����I=�%��ƌ�_Ơ�)j�����\ n�܀9�����1-p�����j"�&��0mL��CM�Dy���R�t$h��WG$�MS3��T�p�Fމ��H���$�h�ZUA�=`-���?$d����O�~�,�"�����e��*��!^Zx�#�����M� ��Î
��{)���R*�������p��r��yZ<�42�;ψ�a���Y�8FswH�]��7g*�7D���zЋ��s��>n�&��?��f��NY� �*�\z��#[�bɕ�p�<��Z5<��my��{����c��2U���Y�ƃD��#�t�tLN�#�AYɫn.㘗�����K��
v����G�����x�7��u�~�'��mx6���i�v��{`p@���7�3�?�t�	$��G s�DwPF��@�k.=��naB�\8�a� y#Ww��V-���"m�D�d��Sk�E�<�� ,͌�^u�e�?��������c�&*�Qn�-]#�o����B�b�k&[�o0P0�Z�ڟQ���k���z�mY@�`�j۵�!ߢ�<v�(��:��)-}r'�Pړ|�����g�lǊl��Q�;!�����@�]��<��3�b���1c�+�!~�kL�@�3Q��_��C �� ���L��VZ �*3��#@.�e��p���B���x�=-���MwmCx�)��

f�$+��b������oXӐ}5�85X�HP}=���|��]T��Z�-�L�	),A9-�j��z�6�7sP^B�TH�@�V�z��A-�O �?U�>���|CN�ø��Ͱ����g���61Q���Z%�g�!�h���Fac�a�*|���R�4T���=> ƽ�_v�t�vP��s�W)����m~wC�7��� 닠��f�ӚP[8�B�g�ޓlﺊ�<`VtuE-�m♆|w�Ǟ+ш��%XV�|�h��QF����z��GZV�`}��a��W�'8e�ɪ�$N◽��i~�����Z��U�,xm��F�O7���*��@|�a�n2����_���\n�YO���Y�kD�!�ؤ�h�6��E6�̗շiAo��(��_�J0]w5�A�G���svl�-?�!v����9�,��I��N�p]Vz�.nmN~���/�#V�qcmh�hb�P����O���5�sK��<�Z+�]���^����h2�.�XMc�u͊,����5X���y���3�"�z�P�k7��i��!����t����K߽"��)��w��afT�G��l�T%r���#CR;�|HBY�Q$�x���6����|�Y�,*�C���,/U0{9J��K9IL��f�V�-��fq�㑷�г���h|�ϒ��W�Wf����q��ԟ��)�Ǩ�	&Х��n�m�ƙ��suYV�؎5�Ɨ�m�F�^�*��F��	�pQ�9L�F�H�	}������x���H�Ԟ)B5�p�Y����1:Մ�1�^/��f�.�ޕYtnM��!��*j/�����|���(of��t/^��ndQ{�5le�y�
�� �0��Y�{��V�+���T�M�Y�77i�N@{͘rd�� 2v���
1a������MܕWV��"�Hq/�1�_�\�ۯo�gB���l���f����*:��8]_;�W����#�'·b��h#u|��K�A��������?~�P��S�^���������	u#�pF�
s+AM��]�>�_.�ڏ�c�*x�����g���*��:
\-& ����?����|�Ʊ��x1%֘�YN� &<�DgN������S�z�2z����!�%>)�'0o{̓S�3�	=��a��=��	ԃ/�%|�C�6ֱ��qb��4���������cL���͖%��
�%O,��a�*�Ṱ:�,��>6w)��qvER9/�0�O�T�7�.V���TA&�=#V�*��M{X�L��Tl�=q��jA�u�&�cN��5��HTI���.�^ο���ߖ�q�D��b���L]�X?��T��CY?�����D<�pIS�pPR��A�x+j�"D���aJsN�u�"�L�5��)B��m�T�%q��Ub�Ҁ�HO]�����,6#�|�����\
���	�_���w���BxⅦ������f���;Zl�6�30e�@�L?�Fŏ��J{0	�n"��D��خn����'�;V�E�F#�Ǆ����݊Gt��^�۽�K�����N�QBoM�Z/�*�A�4������4��-$*�o��&���[��*�1�&���3���RHt`n���O=�
 ���g]uC���a��>E~�:h���zX��@-OU�I��4,x�U �{�wv�!z��qCd|t��kցjպ��f{U��p�����˞'���>Uf���>���'F���� rˍH��	?��.`*��.�Lv��q�@ �w�I�b�;�r=�<7st|Ŝ�b��5����S�~�L�Мj|wB<�����\�塦�ek�q'�R����%�:�#�G|C,�fi�aa\|�o2!e�}#-�A��$�ǲM����97�źc���zջ(������(=����ELE	J�=��\�V��q�q��e)���_嚊/IK�*|��W��^�4��{j�� �q�Y���l��Y,�'4Wj���	i{1TJc���g羒XA�=��`��Vu+<M�:�i�[6	���ˬD�K��"\����A�J*򓗑u������T��
^[`!�~���x�~�gv˗ϼ_�Q���'�c�XnG���=�r��kZ����}����{��@�Jt5D���n.�Ns}�X!*�t|�+9�[�Ͻ� 	R�`<��OI����:���zR�tOkt-= G��8��):���=7�\>�3���FT5t��D��}�y�����Z,�a�^}�(��fO��C���������ɜ~sW��Q��ܞ*�bD��h��m��_�K�� ֖&k���	��.��m�7�*��@�Y�����a[�%�����l���~'�J&)�:I)��#���ݰ��
O�<A�(�����y�M����m�D&�A��$�R��ݭ�
��A<g�zӺ�іw�*�E�����|�̏x�ܲbZ��R�' ��6d�t���i�!*Y���7��x�o(�AO_(��voE;`a��(�$qe&�QB�T����L�w�}�$�X��Q;I\Gm��Ql�}��.�Q�jȧ��:t���}V��x[Dȁ��V��GeߊV���¤��nq�3K�UN��f��Kȷ��Z�	����oi2j)��B)X����}�9!��{��(|M���li�����A#������8�&eki��Tg�5���w���y��VH��*�/r�f�2��.7jor����O�Ik(ح�d�wr[�%*-#���Q鮏O2N����U�[�}�v���>�����/|��p���7a�|��5�����%��TM/�iJmlG</oU����Gюb�!Π��V*If�ɸs��r_|����ŲNaȔ���P�n�A'�Ep�c�z���}����K�F���!tv��vti���?@�.Ė��?h]�Ox��� ���yƹ�;u�-%ʥ���vnZZ_�JAs�tn�{�u�cӎƸ�mk��1�.Rȱe©vh�����ȵ�t����*�����k��m*��{S���L�aY��Ys�wᚵ�ߍ�\[�2.��mD!�,&D
�GP��r���wQ;��^;�N���C3�~s �A/�M��K	��s��q*�2_��f9��t��������6˵z5-�/��1n�CF΄3�{�����
�9�)����W_�<��5cVP����ҿ0#��u�C E��/���a�X�����n⛰C)����1�&x��H�X��^���9�t���_T2�,�@,س_�P�a�!x�HN�&i��4�Vd�&��m�h+�~�]Ĳ�̯�di���b��V����<D8J��Sny�7��A;��dk���=��U�hH23���g�7���i���V��u;��x��.��}:�_/h�p�V\�}!�(�����H��w��0�u�X��n���N���ܔ�0���c2��qi�~�Q�}G^��.��?r����q�@��SN���;�ͅ<�F�Y�mï�z��ѷS ��^��-����U�dHQc��Qȟhh8|`�^~�U?�pjz��]��G��<�ɹqq]��h���@G��ܰa��*Q��\��Fi����b��x�ߐB`aPGY*���z��cvJX^�bs��ܶ�2��W�#*c��k�c�U8ɝ}S1]�i���������3ދ�lw�OG�4P�"
%���#�u��[����X>�pc"N���5����i)A�:6�u�4s �ާO�>&���w�[ӕ���u0�d��<5zԻ��γ�KG�&sл�b�_���:�i��_I��>I���Pc�"����&!�	�R:���}k�.���#}o����/�s���y����Х2}���S��A<m� �<�ӛfv�1�j�y��8J\���m#3�+ϑ�+��_��	�sD���R�a<�ní��`�p��G��(�ۛ���e ��'�õ~�(��l�Z|�h����	ٟ�j1���?bξj����G#��X��e|����{��c"��-A���_CM���.��+�O�8���ִ�x��G�n�)L�XQ����)����(ƈ�ҕ�s��\F�d]�;�n���(���7�P�Q���eЎ&�o(�s���6y�s��\(�N�1>~�$�ܤ�\_�d�i.]02cjHIp��e���T%r[�>
�� ��nS�;�Kh���5������K.:�ȿ�'�f�s�����&d�Ì��M=�$��Eo���K�&�Y������6V>�ޙ�؄�f��?R�����] �$���	y��f�z-D\�� ��9g�D�24����o_n�k{����c�B;�������^��O���R���n�����f@���N�����0i?�G��9>%'�2&-2�@�p��J隮��.�'<~�����GWr��s��ܽ��FwCbA��=[�Z�h��?	�'�%���F�X�@İ�I�a�m�l���)��l�X]K��%��I�8���%�k��/�DMp7Ӵi�c������H�;*��!�vJ��,�N�����{�BO=��0��r���!�?�V"C�jo�^+У�~U���J�'ֿ���W\h�\*�ߤIֶC���	IgpgR���LS���]{ZL ��d�qZ/�D�=�� Jy4����� a[�N����e�����kY�{a��xd>F>3��J�"?�C��� ��`��ܧ$����ӯ'�-8V����������x��b��xyj'��&�JP�źXd�;PYc���Q0���/7k���lջ#��mgŴ&� 1J�����5_�z���²�	��=!�b[��1�-V��K[�_t;L��^�f��� �qV.�c��v�,��W�WvvY��I̠��罉�Q����*����/o.�ǘ�d
�vs�?��D,�V��E��i�wy���P��U#6i�m"��C6d[���]5<	�L�EFu�7�/�sMr����x��6:�j�G�@��*	�q꒒����$!�#�
v��ӷ,It����D!9���3� �u�$�M�s	]�d�ciėڮ�R4�/�h���=�/��ֻ���1bW���{2Q���x8�@W!$�9��j���=���SpȆ��4uu(�X����n`�����ў<W����Cd�x�f^[�s��Z�D�\�,����8�(
�o+�}Kz����ՏG������{`m�·uR�\@��]�+�7�*��7Tg�"^�T�?~�nS�����B���7Q3�걚��긗:�e�p\�禫��ngs��St��=
�x��K��:���V��X�x�!��ϘiH�uzi�Q����������\�5�(�!*i���DÌ�i7�`��_}��W#�g���1Tė⢋q׺��Z���TL��O�Ͷ��u������Ro
E9?	{�01 �l��Ң:�ߒ�������9�T*�$��ô�nd��ag���P+bʚ��P\vh�<�����V^�=��i`��}R��aH4 ���%y8>�ْy��ǚ�,�� ~;
���d�����(\�zV���ԜEwyȋ�����n^;#��tO�d�V�ź#&���o��I��@H�����@ܔ��]���Y��:"P~�v�z��yJ��j���P������f�?�)`'�_���1^��Y|{K�gC�	
$(5T��_��A�y}�Y�L4�(�5�e�Un�S��)	�j6�<G?k�Q��&�G	�b0S��e�E�ۚ�9�r|�~?
�gΗv�ې-}�]j�"�3UE���ˎ^U��`m�C,�҃�"����}�ْ�'��t�k=��6P�#o].�~R�$�
�(uPe��*��(V�d�,Y�m2��y�Y/���g!��8X�s��9H�wJ�c�&c�.[���E�9�P��U�]*�vE��R^u�j�t/��o���\t�[�β�����Ҍ��v��Q�%�{���x�9Cy����_��ni�~Ġ7ۓ��s	�#����ח;+P\�?}e�aB)�T|	sAi��wȝ���/#=n�b#o�8�^��.F�2u�P�:��S[
~.k�-��<��P��{���pJ�u� ���Kgԥ�P�6*��z�}`�[n�=+��KO�֢=�J�J{{ T�Ṅ=got����B�p���2�gL�E0)�>���
-��W���������P��`o���K��\�Dgo&j'���t�L;�%Ђ~�pԈ�J���>w�;�~:o��μ���}����Ɩ��\:��_Z_����`I��j`��AuBS!����k��m=���4�}�38)�Y��w���.8�d�%&X��E��I��]@��A�7����p�
��(����<�T[����lE�̳�`%_}��6OE\ǚ�G�ld�CAab%gĔ�
3�[<>T�'�b�$	��W]i���`W��C�SeN�+H�ҟ�u_(s�S���@����^�]ǫ{S��R>`�a�~�z4�v�w|l�k�(�ͨ�4]���Y���fi���.�ڧ�y�ۄ�]��������@U�H��uEK�'f�p��MMC�)0͛�ɚ,��#�{;�:b���Ҿ������9<�u��< �r��7�q'�)�2B���/��9�A�i#�s�bjhʻ���J��7�S&N���H��^�f�jQ ��遳~=�	�tE�����H�}�HI�t�Y4GV̭n���c� 6�x/a��������9���+Gw�Y:`Y=5W�M��F};�9Z�`��r�;�������Æy��V�W�<��뮄QW��&���܅�R4�T��� ��~�*)W�+�W�[��B��ZK�~��ۢR�<�<n�%�G��3����a��Y�%e`>`�x�c�wc���n�
<�WD���l�)J�Z)�Y�)b�m6jz�ks�<4��a��Sq������*]OY�M�O������B>ܢ��I諴*x���1�c7�|H�_]�@�a���-0�q���m���%�]���\����m��eA�_��כ��AU�~���6��bΑ-o���A����Aہn<�R�,���Y�Ef��I�o��L�=�v�&1P[P!Η������j?�)"��˄���r��o�H��O���Q֫��:��s-�|�! �L �f�����k��W�3���s	����������;���T�4�?L���u1�e�O�����:(�Fo#7��hu~�*�q��@�����j:���YMWl��0�v[i���YQX��I�1kR�P kY�S�Qh(5�X������Ӑ��5��6��2�o4�%�?ts��b�0[ut�S0�N�4d-aV�]c�:�.�� �pʱ�k������MHI�L�0��ل�jO����?<�3��:U�H�n�k"��C�Z��T�G���%\Ћ3�D����=F�9�,��B��b�tWǐ[�V!i�@$�q��Hnas���؉�x(@�YhIќ�a�astk��.�$84e�7Pχ�sx1�}差n��lx���Z>̰t���{�O"�����lR/j3r'Jke�S��E�t��	u��lйO�;�����G5�}PI�|��6���A$�����E��uj�"���_��7��pl�"��$���^Vq��A�_ ����mLû�%	����%� Օ ]����m�d�'��T��r��`��_�gA�xN�b��О���x��c�<ꕱ�޻g���Q��	���8�Yt?�.�<�@�>��cD �/P��ud����I�P�!Bzܥm��"�Y�܇�d�� ���((�mq�'�����^�R'��C��G��B1"�:!O`|M��� %�|���kW�2{����VM��#����e:^')��*���?;'E���c�.����Ly���2!J=�u0�B����H�:Y��:�7���4�>^eK$���mh:��*8�����D�.�)�址��w(SK%9U�&�]� ������3͑,�8J��%��m���& L���8F�K��O]�����|F�3T�;)i�z��� ��W��JW}�P���q�*] �%:v_Ί�/�b��Q=�"+M��g\��'��ꛎ9�:���<��p�r��0t�c���O��-��<l:r.}�X˦sBV1���(�ib'���r���'g�W���o���Ц�Z]��r���g��� ���(4i��uT��3�r�2��p���a��jk�w��j�ý��m#��������L��+|����c�~\����]���j올��x��X(�aZ�v�B�����d;��.���c{ѿyU�i�P-d�E+��f9��=���UL6s���6,�y�6��Y����i9���M-T�[��+Ӊ�ݠ
����5�o�8岧.n}����N�;q���_���Qg��Znֿ��~h��x��oP�"��?>q�(5zT|l�����-�����ġ�V��o�\�$$5��$c�]�¥hY�א/g0D�v�|u.[H"��
d~�UqC��rs�`���-��+,ʣ"y���~�X5B/�J�'{�Ĉn�a�'��l�g�E��.�W�6�;_���f�h�*ֶl��F5�xj�>S�8��@��l��9�IP���L����ٷ�����<ʑ�)K�7E��+tj����d˧���9��Y���hSθr�{��=[��Ѹ�̟~���������)h��]����ù4$����gk�>ԟ%���M�#�\���}ւ7?Z�K��E�*6v�oH�H�4Y��fx�'��{��\G#L�c��+����0*&Q��q]1wO��΀�>��3�
*��e�߂H�����4��1>G$SZD�7p�v}ο����3���a�H�3��_��pe�i�o!=  �]h���{2�R�(F�Q�m���vDC�G��y`e>�E�<��X}���d7��`�~�I�M'3���]�&��PK�	�,� @"��(:����{bw��N�`�h�E�7`h��s2)
������b�V���N��7l<}�����<�J]z���w/e���:ز_��v��s�r����ɳR�WjoǠ6����j�ZW3d�!5��������E�h
���e]��3���Bq>ihT���y� V����Zj[�~�?�����^œ<�D���(��C��bՠ��`�tϼ��LP�S� Jd�������DR������kӾ�gκ\e�q� �,gE�)}�Bn�r�gn�1�D<K"��Y3`� sç��#�����2���hS����6��1 ��*���b#�*�#H�q���_N�2 �,n{���G�l�[f����X!!D��	����?�3I��������3HsBCЛE�l�HY�V���Թ��JQ��Jb:���)�[���2S����g�eW:H~�D���)�r�VW!�@�-�L� ���ƸI	�ePq�
�h6Q���p��ۻ�f�9,-�"���Ѯ�Wu�J09���t2��p��k(����r��-+J�N� Wn��#�A��*�q��)?��lm���j̓�
����
�Tm=! �y��?������d�f�2_j����+&�l�!~�A����	�P��w-�6Y�{"��u$V-�ċ������b�*��[|!���>8�z�d3�=���)�&`� ~���d�E1^���z#�] �~7��$Q��:]/7��)��I��8���2��@$���0��j�O��z��>���;���Q��"X�_6�ٹ��n��m�#̟�ϳ#����?�MBT��T�����H?�,�����s��(��s�m{;���\��z]��Z�欀�IB�|�����i�%s�ˀ*���w@YR�p1��­��2��*P��E�3���xJX2�x��/�BYӢx��̠�%��y�Y)վ��HI��]%a'��oC�Kd?|��ʦ4���PaK�Apt�V�-��pt�w�^�����tE�^�[�ŀ�7@N��i��+�ʌ
$�Y����ŕ����m&��^�#o:uY���5�o�{]�� �O�Ԝ 
�d]�;�'[v��h���4'o�q���\T��@i��S������r� ˰=���X����r��`_�C�iE}#￶��� �`۷ﱪ�d1��P�����::��FC�8�9a���æ�ku{*aMyL2��@c�CN0�)�)�� &�����vs>��R�h0�������c~��I[��bƶ�9L�V���)���]W�ˉ�"U7�1�=àp;0����
|�=y\ߚ�mW��41(��oID��u�����g9V0�@27�fs{j��ջn�ώ<�A�$a�e+_�������� �D���Y�d��S��+iɫ	<M�R�sv��^�M�݉TӮRJ\��j=<�J&�J�����n�zݫL�&�tL��I�F6���3��7p^��W��N�eS����I���iƆd��"�n�M�t��
�P���jb]@ m�} ���E�����F���%���#.����~C{��[!���V��)=�����YG���&�9�~zi�թ�0��|2��Ɓ�s1M��GD�x@�������[�g�V�>}�K��+�3��Ј�H3�E댿,~�8���6��_���-+{4�L�yj��_�:$nuzh��������\�V�l4�-e�{]��Čq��Ub�8�`�Xj�**aBH���uT��?�Ĵ�E&���#-��&|�?>x���9q��5ʢYK~?���F�g-%����s�rjF����(��1��mv�2X�q~N�����wt}�����N^���%w���z5ϭkaS4�����w��(u�u~w�)�*�����mH\�~z&)K����-�xZ":ܢ��!YZIU�@�lng�4z܁W��?Z�����~Щ���;aC���_J.�<5��=�S ���o�Ō��x @Mú��$�-�,&�".�gj)6����,���E��xq�� ]W{���0�s� ��xb�@�#��}�oiD�)@���b:_�ҿ�j��3�R��e�=��!�}�����Y�<-n�0cB�w�f�x��S,��ּ�˞,�p���C�	a,�d}-#ճj�I�P>Tu�U�+�걷�5�Kk�^D�a��Z�"�'BQ�rK��ͯ��0&���{�8���,a"� �������E�𚷖�w��_�\����;xl6l�Y;�0
L�����ˁ�L.^X�#�9X<r��5���L���TݙbA�ٔ�hع�Aٵ(6���y����AvTT�Ȫ	��<"}�� t��YP��m���Z�8SS���FY���%�G0ԡ9t}2��]
]�
��*�D&�Q�w6F�Yg�P�s㾧_� @�?��1���Yk��nZ�nJ�üծf��������IL,��M���T1����J�,��a���2)zX��z�oZ���
�G�s��J�#>]l���z����ڼ��b����ڻI��D�-8���*�!��&(o�>S_$ҹ�
��oNx��ҹ�+Ű��I�|�&n�%�Z��O���:�aИ߯��$��6O���2��	�{���Cu�=F�x�*��eh�+f���D�ˢGE|�,�����>�����j��Z"m���S�d�ɿ%T���y�*�vؐ���,�)��?CӪ�ZHb` |�P�O�m����MWB���_X���V����b�_Y�D�ͩ��y�X��t0/� �w�	��hG�DL������[u�Ų�ʻ��0�eʷ�\��JPC��J8�Y������`���xD��ag��*����o�5�n�����M�l%��UC�F3��L�K�P��NYSz�8���M��[7�8�O�b��g�^���W�7�[�����"��P�*�/����å���+�M$ox�ײOYt�q�O���m�\���0i��؃�<JX w����M�Q1��.2���3ץ��y"�^i�(�5Ygf!Y{���S!�JN��c��@W+,�?9��;{��$Nc���=��u���ݛ��`c	)F�ɬ%�\��@  ,q��g*����q���b���r�t(.V�Օ�g�#0d<ESk��{__�'�~���?� ,�_2OM9�p.�3���v{1	*��T��BGXc���6CB��>iZ`��>���K���	A3��0�g�p���|=L�4�Ƽ�q �B��s8�F!���55���6���{�:@ˏdl����(�i���<��Z�Ueuz���#q�
ͱXB�ϥQ6�����v!��6�]��:�;(ׯ?zx[v�!"�sp��zH.豦"�%d�-����/���FR�UY�~U;=� rG�7���b�9�v!�Q$YL�vz���	�n8��Z���X����K�$�񜥁�����gϣt�eH��w�t��G�P��ӥA�������6
c�5�hh𳃜�b�3y�
<���U?.��q�7�.6�Ư!b.?����M�<b��1�ab��h2]ZZfs΍,{�3`����[����o�60��t����J-f.d�.���t�=�Q��c#"�|fP`��[+����Ý�-�p����������;fq#Jt-��)�!:-����p,GE�aD�߷�1�ǭv�H1�=u��̨�o=�q�곽���\x�/���q���S� E��]�4$u5ɟ�g��4���X@�Zf��R�i���:�=Vt&�D�2�M��L�iL\���*=0�&7&�15`ۺҢ7��7����)
����]��0;Q�&n.���d1D� �(!:v@���h�<ͻ�!D��U]�u�3b��g�?R&�&F��֍rK���2��rC4TېW��g�+6�2ȲQ#���k N���ɹ8�j�
�VZ�\}����9q��и�G��ݪ%������qezE���R@�8�(���x�n"
��7�[�]-"f� F��2��r,gJ����.�n7�Ʒ/rQ7;l���}�����t.v�ja=Cʰ��H`�Ϗ<�5�A��aV��ʰ5���rD���ۆ�*��#��g�΃�
.�e����#j��C�������|����<U��"��i �ؽ���/���Y̟~�'�[q�[Lj��B���z����h7�(jH�s�־2�j�����Kh비�ݙ��1~���)B/\�md�wS�׎?���?qr�T#&O�4o�o�&��n�;g�Ȁ?���=S�wX����9�D��)e�^����\.�6�	G�Oͨ���y(:#1z��˝^�q�_�imM�3�&D"�'�]<�t�;Ag��h@�Z�'��"k����Ъ�q2�1�r����*�ݗ2ߕWy��4�~�J��t�ϯ�hN%�(o���k��m�\r=�hY��@��9�v Ο���F���6�?�ܽ�H��<N�~AmS��p�?�Mq���Q�Ɛ؅�xQ�����~�V�ݗ)�\f��e�k6�D�3&����y�-�8����i��*3J��OB!���K�c�`L2u$�Ɠ��Wj�^?���}�LQ,�� ["N�N�װGM�6;���G�$,2e���'���|�9�H[�o��1��!g�y�i(]yQ��]�h �Qu�L���/O�2�yR�>[�b�Q(i	�t�^�����zTme ��X�����m�]p9p��ć��kˍIҎ6-öOGl�x�ؗ�juE�;�K���oe��:���V�Q3�϶wR��q��I������;y�F����{ۍV�C��"�M�{����Z���ֱ�SꀹÜ����_-�ފ� ����?=���b��	�It�;�����e�͙��JxQ�K1� �-��!�h���1�|1�'(���̦�y��!�}N��׍�9ˎQ;96���
u�jv��.�@�997��`�K��7��/=���H�'rxCð�O�%�����w"	�u�=1��*���Ƽ���W����'�^�j�揂�ʗ�E�-��Ju-B�`�
��y�_Ǥ9�cEd(_˥A8}�5Ƈ*R��X=��,�`
 �����	���J����f�A=���Λ_y6bR�|��wt��"�a>Kp;wJ
@rU�R�Zq�&ip����*&�բ۝�B@~�p�a2�/1�Eͩ���r�s�����5&��^:J}��I�`���Rjr�^�	!V~�b���܆��[�Q6VR��+��}���-� S���`XY_�2<��E@/$t�9��ذ���|�g*�3 ���_r�	��8o�XH�J^X�񱚜l��u%*p}}�_J\��F�:+~�4_�<ͻ7$7�4����g�%Q�bE�n�Oò^K����]y>�=�oL��b�r�yBC��p)��:�B��}w�;��/<��qоs2L��(\'�(��8܏���ek��:� 9���h������J�e��V��R���y�#��ڱ�3���b3.�.��U(�1�/���ʦp��@�=B�r��u̦Vǂ�,�y F��C�	�h�5�_�t��B��a�C1F:>n����=�[3����:�A0e�`��wn9s���s)��r��b�ˬ<����p9���M4�k}�8�9�ϣ���>x6a5W���&~�<f��g�{�s�I�/10����!�� {��o�ي���4�"Pc�(�}\�tjSϽ�|lCp*'����,M��>荜�qM�M,� �Bb�7n�,&�4j�^��*v�^��ǵ��J��t�+�{4:>q՗ɤ)C�#��#*�Y�����qG_B��jŪh"J<ekYzՇd��J���c�����	:!���0���J�:�U5�h�8Y$E�Ѭ#�-������5��6B�(���t�0A,i�~��'�=D"��g"E��[�3�.���A�Y�P�\
f8,ʡ>��T��ɭyi3k)GZ��&`m�>�F?�Ċn����D�d:ع���NT=���������AI�(���C��뽦�qx>��,�B����w?#���&\:!,���)������ی@�N ��8^���b
��hz�Z6F�z�]�Z}���p<V��ާ��~�5v����kX�fHd��s$�<=���FDę�|�T1�*�I���6e�A��/~��[k�i�&|)K�m�:��~�!���+B_�Xm�.��B���{��C��_/�̟�%1�c�jq�� ��Q��||ز�#<b#�w����a���z"��w���q-q!i��ٙ4>�V`~�i��dL�;�e�ۀ�m�?���EJ(m�v\��3���1���c�;��4C=6��!F��NH���Y[�\Mi��N�-{ma4{2��Q���t%�0���~���),Ѡ϶��t�4)>^*�uO�?�Ƚ�n6a5�XMl� �K�X�2�b&s�����7��P�I
����bT	��#"1�i(j��a����ksc66`C�� 0:�f�����SR*��O���=�c-G��D�8m���6op%O�.�vl+,���'+=�#~�=�5�$�ۏ䙰��l6���p��EX�
���Ԇ�8#�p�?�o�������U��΍��;���in��r1 "U�}�Z;��he\�i-]!pL�f��z�og06;��L��1�lY$x��������ZU��3@�����k,�*���.`f�X*��I���X�^���mK)��E�w��k�aG�{� aM�����E�eG�1=���ڕ�(�꺂4/�sv��iH��J���U)o�CT��a�̿y�Κ����EOW ��lؖ��cA?� 5W-����9�ý�UZ�퀆��g3=��w�� �?o�_0E�j�D�:E�J@��?.�R��|0n ��ˈ��#ɟW'��ǽԲ��B�y(L������;�����q�����8�R�O�9��~���7/jBr��^���S#F�>f�?M�W@�L�\���U��Z�>e�+��{"^⾮<��K����D��y�2�]B�8��S�ޭ|3��q��d�$,�P�|�!�=��9�gR�]�ܸ�.�8��UM��X>���TG���b{��ڎ���f�h"�R���D+~v��F"&�@���M���n?r�eɖ�nI����Q.��
f��Nl�~f���i�4r��M2��U#v~�aPc�ɹ��W����B�N��9��G�qLo���h@�Dv��C��E�k����������Q�o���:+0^��Q�$]�.�p/������m�JA�p@�m����6|&n�e��+èn�K������ry3>GW~HU��%�Ap@'���3�?�&���N�ۅ�'�$}��5c:�M����t��I���N���d"�ʷ���pA�RRٛ���0F��S9��W=$OV��r��fJ]<F���D�q�u��O+��d��_L��`p�2h�OS�����!��XQ�(���J��4׃� �Sہt��o*��1ج���w��a4Q��fք#��NУYG�Ĵ�`�#�#r�V�P�1\���xϲ~Sb��שS��	���͗B���o�'�uE��ч��ӱ���%�[5B�b0ͅ��xZ�O:����c{������/�~?�a�	���iL���!��4���=�B�d���G®k�Gw&����m���V{��1p�e�����䇃�	 *�8�˹�DAtV���b��+�S��u��l<�E����6վ䘴�ڊ��"�wQb�	6�b�Z2�u	�K�d�ޯ)��(Z|SU�{�s��m=W��� �"`A6d5؆A}ؙ_)�y@�L�`L�?]�="6}�`OY�Q�)-ʹN�x-e�	jh[�N� ��/��]�?�i��\:96#g����ޤ���>K�F�^`�rK�P�a�M��\>���$��yL<��A3HRg�����_�V\F��g����]v8�<��mj���2����&j�Fƛ ;�FP�-Y�s��B��:S��+Z�/<A�e�rǠ2	��rT�?���%,3q��ә9�!}S�R�-}-�߂�Zju�����݅�h*�`�Dr�&�ῈVp�����s��n�h����c�+Ck��Waᎉ"���!z9�S[a�0E��ٹ�ꖠ+e=fG��@�B\�]p�*pAR�����>���zL@V��o��Ѹ�h/�mO��'[��]_��w�&����1J�2�3#ip�����aG��`�1^�~i��it�s�R�r:7c�m���b0�!f�
���uT(DE�h� :J���g�E����W�&�����bH����<+�7�ru&Eyy��=�^�DB^j����'�Eٰ�4��IV��3q��{Φ��M 4�F�I�J':�`]��8n��A��r���n<��å�]��AagR�o�)��L�|���o2�����
�7!�&Q��bs��C`�z��*����4"��p�(6e<��T��Kԕ{��,e�L�s$\b,FB�D�J��fMu�]�<BJ�P���\���X{����B�r;οT�'�wu�-_*���T�2�� ����W��BB�̈́���ޜW�FI���t���KPS���2�3thy\	�~�8Q��zVn���7��C˻��+RY$�>i��>k<ש�Y���>�%	<��aW�6�K�㟨�2�F?4�!�N-jU;��"t��]�Dף����w�+�#�Kb�k���j?r���V�]��In ���Ai��HQXU�5Z!�_?�x�[m��y�H�z<Y����Nm|.f���.�?%��̇ky`����Xގ˹��E߯|�b8%���r�Qd�E�K'�E�ܱlO��C�ޗ��	!/6��ߏ,o��]d�x8ت�3F?�y~��C/�Ԍ_��2"�4�]I�0u���� ��e�0����Ǯ	��6
nW(�����`�^%�������S��G���M �ǈ��$71W��'�nmop^��آ:`*2/�����	z��Q_� �j0v�!ڔ���D!��X�7l|���� Suaڇ���6��x�v^�LƎ�f�d@���	�t�:ҥR��p���u�ͼ��M�	�;���A���u����J�&�Og��v_+���L��=r	ZXh�@��֡6�Å[���h�b@�"ʴ�M4w���X&<��ⲗ1���d��y;hXD뚜V��A�L��ڑ�g��MR��F����������=8$�\v�5R���o�h�o1�I܊��!O��/���Y,�>ʚ��wF�	8�9�r���D�1?���/��Ŷ��3��Ds9da��~�d�y.SC�~C�����'�"6��i�{���>��.D��T����N����th��'��:ϝ�2���56�:��MҤ��RN�1� 
�>���06z��N�	c�1�pdl��_������	�z����30�I�m}�+V��{�Uw�R����E��d���ŪV$W/���x��V)�#u��`C����2)VP��01c�h��ʤ�H�AlR�0y��o��r�q�%���*�&�Zm���-��"R��2����K$�UK�|5,鍸m!Y ��
�� ���"�e�21��j�_;�>��&HE�a$nx�Ң~;Ey���r*V��L�n��O{2;�w��*I�_�IY� ����
��TP8I�0�|((��$�f�؁�
����Đy�3BE..�:k��Ա4���	��a�֧6��\؈���!�3�9�<_�	�sk�*��qE2��
�cE��w>D:}��ҷ�2�xr��7F���"�X�olJ�R��vpΒ��6�h�IP��ח��ڼ���a�_6B��N�ѝ�E��2�T3�cnٷ��n<1u��Z\So�߿G0ې��Q�{T�}���C����e��4@	NH~�\��Z���ߎE����B�Ψe��!8�X`2Ka����=��w�'6:�@�E/�V�z^���Q�=�����;��+=h���бo���J��h�jU�{�����I��*�*Ὸ=nMT�:�#�4�vp�Q��o���5_���D�f�ٚY�Y�Ñ����|�B�cm<�Pɲ��s �T4�.������m���`�g�|p "���-檯�;�?gKz�w���8w���E ����B�4��L�1��]�p��$�F�� ��I��@8x����@l��	y���*��:l�+��q���(��B��{��
c@jFlh[e�o�S�B��Ow L^���V}�5^U�+�Jw�bu9>�b�|(���^��`٢�R7Z��on�n�Xi-u��89.碯B�y�tڝ�߅�x��N�N}��"bErc�����R	��pzr�>�4�!툏�Ai�yY�L�� �D�`oZ����"Z��!� Hk�� u�t��J} ���,�@�0���2��Z��SX{ԁw�!L�=�����eYqͯġ�����9�͖挛��#|P�J�x��\�Ǡ�w��c�/K��]�"}#Y�Bd����`�Lm�� xi<�� �>�M%���.{4��������Ѝ�g^;���ڼ�E>#]J���^.�
t��r_[�k��\�P�5�3���P6������V��/��h�g�
�T���aT�b�߅nC�P�ȍb',T!4�R�d*��V���]ڂ���uO7�0��yۦ��2�R���,�/������j�*���"��NEA$ hy�<
����b�*�i�pp1�- �2���\E9����F��P�e�־D����^@����I�!�5�e޷�^�����,#�����S����XL�y�q��������Zꕔ���X�RX����&T�Q����&���$#�0��i=æmV���Dw���	SdB+ߎ!��t6��t���+�H��yfB����n�������n�+vঢ�f��瞫�Y�I_�ͅ+�� �_��	N�\�v;���n�ϼ�D��r����{j�Y|a�11 9S�t_�Z�������+xU{m��"��*9���M(����j{%I߁���q�]�םzZ5gzs1����_�ft�\ 	�a��H�:�~Hc̭�Э�6�x�k��H��=l��k˿�m�����
p6Ù���GeX��̴��V�b>r�HY�nע�����%a:�#oۨV��g��TrE��}��-P�'�&��S��� E�1��_�À�b<�t2�Y�E��<�	�;`Jd �+r��^�C�\�/wy��-�/�}"_^H���ƴ��U�0}yq[@������)t2߮��Q�����z:R?h1�V�����s%�r��O��z`C��/���E��/P��
c��x���TK�
/�TX��Ej�#�yխ���]�nc�0�����؜���C"	�����T�����6�k/�LA�ńQ�?i��}�Q�i[/RЋ-τY ��g^�)^ױR`:'��'��5�Y������VE:K$�C���Rx$Um�X`����A�?�rS�hG��I0V�_!%\��]�N��2��eX!o?������~�ls1���ϧI����e2(�HN9��;f]��1v-~�:fԀ��=^K';1-���ݒ�J��a�%y$�5�Ok���^jg�ˈSӤ�",�Y�tOk�oTj	�i�s�p�M�
7 r=qq�"/;�{1����@(O��;�$��i';�Ovⱙ���[`�&��!���d�ť�]0�cpv�D���h*l�$��#n�{4�&g���1�^p�!2A�V7 F5��{t6.���y�16����K4�����-�l�vJoPԅ]3�sz�#��$�z��Φ�'����M�`v�O��Sժ�?z��r��I+̻�F7?�>�p���T�e��1@��[=*�mO��`?M�'=$`�ËƐ��6�pty�� :. �IRQ�%~M�[4J�.�O珪x�6c��'d�O�����͖��	o��OV�0�=����zC���9�y<'n��h?� %���O`o#�����
=���������֚��r1=��z���;g��c ��\�@�P˦&�� �㽲�����Gto����(�K�{�Y��
�I�H�'�Z���R��-دh��l��옵&Gt��<36=���LJ��M�Zl��[�oIA�y u���V�_�p ��^�D[�C��%��q�Į�S��W�<�%��:���L>�K�r j����j�7�k++�򌁽�	nU�$�˙���^`O�[��1B߿+���?��12��� Y� ��$�;��\��V�1�Urlu�]&a �����j�K�q�O�Q�7m�B��ڻ������'��fl^R���e�Y+��x���{DL��Ѱ���e�i\���MV�;s.���2��ۜ�'s���tb"���}���1�t˪���cتȕP#{w5Ю����0?	-I*J�3�Y������`c�ǰ��M�Y(�r�ڥ�ƌ��YC�&��o�}�C��ra��5�����+tM�׫CSh� 5g>GwB�r��ڄ=6�bQ��s+�װ���do�3�^Cj�� c'�D\��|�hCmഥ`ܩI�ePȞ�����56�����4Өݖb'0T��:H���y��)�r��f�f3�����n�{�z}��6ѓ_ܫ��C�g#ժ�^#�T����Ӄ�y������ ��ZX�c��+
�"_�I�T��O9W���B�F�?�o��;�0`Wҕ�[����/�J��d!!��i�_�A( ����7�`ؽ��2�Dg�n��/����~@�D�T�_NEQ�?�@%^DD#�1��K_g١��O��;#V+SF�Jd����~揑�AQ�P�GM������L$�2>ꈓm�������a�pɪ�"Z�{�6��B7/�r7)���ګ�Ff�H������2u��d�AK�{T!ƿ dk���Ta�ˈ��$��NH��2�Rk���4�&#��ֆI(���O��D��+e�r�7�s�tQƘX�/�	��J5�B-�!�����G��`�Z
���w=��:_鉘�C hm1�N��܇��oӠ����RI�5�Vl �b���t$ׁoP˪�p�//U��j0�n,M&�lt|h Q:x�*���4-��ZlЄO�a��G1��5%���Cc���ѯ�V�z̙(}����0���~B:��Hy�'�s`�Q|�>�B2H�s!pn�:و�'��v�V�ۮ�A���[w2X �*^�#�Y�|�T����Ѯ(Ů��Ā���*��:a�~GM(�a��FY�����F�c2#��߰������7����j���Y�
3ep檲I��E�2�q�,6N��C������{��1a�g��|�Bt�0�`�ު������$�o��_�2B����ŧ]��m+�R��,S*\mŚ#�a���:gMw�䷄}��U���{�(���h�ƕ�����3�)xXR�zR�ŷ��:�6M�P��]�X��nq�Ve2���z�?��\8����_EG� ���	1E��U#�)]��M�	9�i@��o��Gj/Q���̐�0C 4��v����6���%Do#�$Ot����U�Çd��*�ꆀ���@b��;�c��LKm��Os� g ��JH�a^�`�
�Æ!������c���@�[CٰZY1xma�>��
�&��������T�S�B}jX��W�� ꛈҢ�l��uxc6�Q����ֱ���Z���_��7��5I����#+�1�l�f ��L�R����צT�*	�sC���vU����1��k�ʽ�-m`Z��Pդ褊DL�1��SAyE��,+�¯s����:��d�@M��o��Z+��@bH �G�������Ke�h���@wf�NѢ˩����Wͼ $R�O�$O,ŏ���ޒ���0���rӠ��%��qӡr�o��s��{��L?�����M=묽��2+��&��I<����lC��U&�A%F>KC��>x#���5�Dș}F㟔�"rwx�ۓt���@{�a��FJ�|4¹N2�h%M���~*���|�%>����u�+��&���=�?���5��#׾�U��x�_$7�p}�<\�WP�i��a��"+�A���T)=)u�!�Ľ�/~�g|���?NѢ!��(����$�p`�[�PǢ�����i�~��K��u��T�B X�ǘ�W�m�g���qזt�@�F2���?miM�y�3ϳn�7=]�<��)�6h����?
�^Nl"�=}t/��$���0���X a"���*t�9�'�J6��R�S�oq�7�@WB�l f�$Ae�[�1�9�G�/�g��J��'�B%�hc����������J�;����KI\!���M=�DU��Nd��f��)��i,�1@��@�7m��/lt�(�{���r��]�c���C�&w�J����m.�}�[]��7�5?�u�/�oo�43�9|n��(YL¼G�)*�E?cя�o0��yU9�NyY����t��ܠ�ut�h�o�Yb��9O�h(4��]M3S�	��!�-~�l��^�~I�$q�L}�8"��U�:n�v�m�J��tPp\ϰcb�D�ʪ�%��B8^��`t�c�6%���I��m.��ᵥ�!���� ��ء�1��� G���BѡZw�s��4�o��5xS|jH�n;��ё�#�I�����O�R�S|߉
��9|�&T���'YX��h��:��pk����g�
���0������x��^IZ���9"U�����">�|��{g�h�a9z�~Un��u���z�6t}t�9P���7��?}|�vo�J���(nhU�>)�v������nGgֻ��(O>y�O(H8m%f�\���v������lѸ;�"�� |���u�����~��܋KW]zc�SR�'LO��۳�U��n�Lk�Y��ʵGC�H��u�B��FP
�%d�_[9��0ϳ��.�&v2Vo]���Vc�>X�V(�V�X.+LX	�����](�h�S>�)�E7�71Vb6�������J���FWR�:@�4���P|q�8&��	��KU	����Vh�ٔ���;��߭�6�!8'7�	��p��H&�p[MҲ�2�K�qͧ�/�}�����K,�lt'�d�l��g;����9����j���ʃ�'A��e��n폂f���(׺�P�B�qi�{0�B�k[��{�?E�\�����,�����;����_� �j���1<ve�)��5�a���e4Յ��(��4��w��d�V'�T�K� vn�}�r4	$(S'LZSʈ��ba��R����cHN�۴�8 ��V�L���7t��7_��2�'��=��-��gk��e��	�~�-�̟J6������I�R����Ɯo�Ң��[�Iqb�r����B����f�����_Nڞ�KA ������%tL�3}8�mA7F#��y�Oh�3'�G&�t�4���� =�" "��_o���7��w~��}N�!��د7�J6g��gt6�0g��7}o�WF��v�Cen��ni�NuF��T%4�)�s���i�kt���)����P�`q���`v�+�z/'���q/�P�+��^�t��#�縗wIj�>�6�V-����
��k���iw���gg�9f�}�ec��"W;��we�j�./⌄|�:�^��yQ̯��'����n1�^GZ��9��BЁz�>|4	�H�6a��f_�nw� � ��!��.6��W<����n����|�
.3�R���P�2�s�/�w������5�ұn���)���Dri�J��SB�(�!
�dX��ceN�M�r/>]��ȍ+�2�e�y��Ҷ���B2�W�Ä�X�l�ouݥ`+���9Ϸx�VAN���*��ق�{�����,�@/�+�_����L����0"���Z�ozw�]��ݐs�����W��Ν��T��n|��2�8�Otá�Fu��S�!=&`�h���~]n1�zd��f���kwy��K�����]��9�ҹA�,��ݿ���B��Kސ%���Гƽ��K��J�|��"5s��0Upwm5yf�,�dfD�cH�.�Dڃ�H�����&�=�p�����������97�M�Qz�����67Bɪ"��q�iPw�2�u���4���	�icb�9iJ>mh��b/j�����8n���P���%<eq�lʋ?��G������ �ǋ�AT8���ҿo�^b�w�f?����.WĂ>�޿_���NU,eX�i�-�?�(��䜘x�N+u��[;&v�=��9%����4|�*��мg�(4�´���A%�Rkw�	��^���	Vܸ�[�
�DѤӥ�����&A������ZDXp�M���X7��Zs	b��U�P�b�6��S�ea�@$d�C7��ϛ�����(pKPF��*�Q������2����_��/�S�>��y�H�br�zWҧR��$�+�G�,[�<Mq�f��#
��f�*��+����9y����V�D��g~��*E�'4�9@��Ԥ*�A��ťl�"���BAk���᛽���i�͟S%3D�J�g�b�:�Cu�=^Z�������,���E^���<e+&���hI�nD�#4*j��Q��F{pO��Şag����e� �J�_����&�"!�S�He�n�8GlQ�ng_�᳔�r=1޳N�i����+]2�m	�7⃾3�:�7o#~l*U�H
����P����hj^�G�{}����u1����$��.�g�92�g����c��n�|&�~��5�;qpB&�� �6F�G��V�nڊ��Ȯ3��^3~��Ter7<njڽ�����E�o��z��?�8v_���v��V�C·匾���J��`��*K�l����׺
!��mfp��a�]}�I�;��Q2����׌�<�=��]nh��.j�"�zW`�X�_��R~,2~�N��h7��I�wT��n��{��Ò�}���"Q��
{I�ԃ�b���:/w�J׾��0Mc��f\މ���^7����I���D�pc�q^�}�5�\�X�+�!w;>�� ����=��'�$mQ<���Ύ��k���egn
���/@#t��S��*�-�_�"׍D�}]�?���K�um��n�/��n�҆f�W�������������&2�1�t�<�2d��)���B�f� NCϹ��"���cO�9g`1��,,���bX5}:��cd�(��F�������7���l��Ж-,�Zy�g����ܡ��$�9�h�}�u|�_� �	o����V�`����(��}R�՗g����z� �(.v�;���" `͐h���;���Ɓ��Ũ���ʨ_���>���잔�ȉ���f�92��#����'���j�WNbt$hd{������
��Ł��0�}�,pvk�m �6��UJ��غ�4��R�Zxf8-�Ϩ�g����z&n�R��c\nN%��|���\ ܢ�?v���j��� �O��*�'�W�G�ӈq�hr�9t����D��0������4;�K��V�+��e��pXsI��ק�Q$ڝs��1~Z!�Gg���0>Kܬ\?8c��3�7�Z�?�AY�����<���>?���	����<�22=��ɏ$l�����iK{2�@<��>W�+JD�J+���!.��Ck䫐�Ba�Gn��q�<����`D����\��~��Iא]��=�ں�C�29 +��%�^Jr��!�-kO8G�A��X��͌��ύJp���n��C��|RQ�Ӛa`��T���u��j7�Bmky�\;D��A����-PkE�axX�&�J`�qS�L�\֍�8L�)bR�}M�\���vt�A�ss53����x�D�0H�� s��[�x�&c��c�����F10+��g����*@b�hjT����g(���,���w�(oZ2#TXn`�c�G����i(A�s��	3xfϲ�Ȅӑ���P�O4`�#=� }�K������e�r����2Id�����2o�|s��sv���ܒc�Rg��Z;m�����DK����:�!%�q�!�D�BqX|jho��� Lb�Q�o��g�����.C8�;��B�&Q���L+��T:�����;��P-a��H+% Amô�9g��}z�������HG'c�v2�"��\�<���{	����Tm�bƮ\��lʑc��I���
?!�~mP==$κ���&@NX�#g/���@����芍�k�)��mt���$�����F�]�
H��Z0T��,���i2|���R-�W��/5��쳹L�朂	đ��ڻ�*����f7��O��l�%��u&;έʉb�.�fE];�`U�C�7�������`�AԤDeqZQ��ǁ��L'��I(� �6ھt}�@������S�v}F�l{�3C,e�.x ������8������r�1vZ���L@h}T�q9˻_n�<�jb�ƌ鷥�r��-�V.�39�Ug'&r+;�$�Q�پ%J2�{%`_�a
��| �\�[��h�/�1~/�nV���5�_��&�3�(���X[�k~�K:�!-�r0�b�rM���Ĺ��p6�̗:��.�6� v$G }���D5�>�o��3��$�2��8�\��~|W��\��/��u����*�s��+߉���Mح"�< W]�(�p��#O����P����C��;�UXW�X_>�������G��DM
������9	����;����tlݙddQ���q����H�/�"yA�lyBVX�O~��@�ɍ�TY�[ȉN����I��93k�NN��nq� ��~�!�w�o�!���#>�@h��k�hYBd4����r��%M��߼k�J�մF��ϳ��x$ߖ� �iq�<���2(1�q�Ip[c#xP(ʤ���d���s��?L�y#��k�;�W':�r���;�!z�d��yJQ����P�6�[O7<\�;�<�w!��ZLg=���	�Q�coq	�^m1�R���ރ��8�c��r���+s!>��
S��n-=���Soب]p�<}�'����
�\Ѧ��f��	���)��)l:G�-��Ǿ;�Nj�\��-�U�������^���![6����i�nQf��GfF����zh���G�ֈF�5�g'��ޯ)�˩ĥܩy,��F�f٘�b-&�} ��`�TT=2s�JV|��a<�Q�n�Wp��JJ+� ���
OVO��v����X��s��L<?ȄyWי��b�-��X�۬xq�ׇ"*��H�*2s��αZ�tyd~:VcQ�+�YjJ���{}8���/V"�S���*e���Y��W�����۠�,�����9ጢj���%�sҰ��蘟~�·��%�yBc���S��t��զ�kdGS�3�̘>y�����g��i@�b����9,)�T�Ew-H�j�K�Trx�P�����������H�U����X��EF��(B����f"nҲ@�A�9�Re��\�(m%l
\Y��'��U�Lt$��k�QxK��Խ�A?vO\��i�i�mGȦ��(O�&Zkc1>3*�F�#��e�]���.��*b������YK#�����~��C�y�QL�*3���rU@8
���_f�`f��l�tX~�z��� %�
P�8�e��v�#tZ��7��k]�}�t����;����T�~���&���Swa$H�#2|�[�F8H�"ۓ3�ސK�c�&�o��_�QU�A����ʉ���"��G\^���>��:�ُ�cK��Y�g]d�Z�J �f:�L�`J����y�ȱ�- �d;/ǌdv�k�ŀW��3=��}���[d�����w��+Zt:�.�ìm��
6bT@o�f��~x�z��ʣiK�!��\�:9���$9��y�� ?&[(���/�!��6�@����A�f�и[w� ���AI-��/����SOS����P���E�F���c���^��
% ��޾�gM��|����ZM�n�%QPa�ښ���������e��%]8���[8��vy!���3^#>ʕm]Rz&`|��A���S���Ј��F�x�����1�;S��h�������T�t�rQ�Y��C<�+�?�)\=��8�au����m�DoP>�'�3!g9��tnK͖��Fށ�1F�
��j ��{̣�/��@$fB����@P�)5\�B���L^��n� �t���dw�����r+椊S�`8Q?���6�8�[�4=}"��/d��C�������l)�" ��>�(vLm�_�2E�=����"��Bm�hQ)CqՊ�ۘ�|-�����\O�@<I�;��%nҽ��E�$�c,�����=��]�������:)Ip�I��vu���Y�Oήe��v���s�a9�����eM��ʵE$O��ku�2�'/L��knǭ0]�ǫ��u�~࠙��~(|����#>M�c`w���#��&�k��\�"+��;:^rP�h60EA>������x�3�f�8�, f��3>���B��.�ރ-��-�nF>�y�ʚXj~�;m������u��gTM�a�9���5�@�tx�����☄<�2f�sQ��Y�<Sm-y�o�/n�{IÀ�o/�g��nA�6K�ζd�������i��v4/��������u��ΊF����1�N�F��(��+����6��aF�Xwp���k-,�Gf/ۭs/Ō�Y��w+��UAA�y�y.�z��qy�4=�+��6
��K�>G��>9<b������7d:�I��^jV�]V��$X9� 0hCM�
jv4w���_�����a/����`k�b�/'&�,�̨U�r��ۡ��Nt��sŻ��!6�1L�\����D��Đ�R�&��\��X��s��Nm�#��0>�ܦ>��7�]u>r����IZ5�1rj)!��b�w�(g��)��,G5澊E��j:��3&��m���E#U����@ŗҲl�l����MT�r)��]&N�JP���V���N���nY��F��><.��G�����0�3Q9 g~P��=Ⱥ~��fK�P#=��l�ʮJ8l�>�WB�/���ۚ���"������V
鍙� ]tԷgT�h��k		4ɀy&��3!�܆��#����Ý�7�B�����Y�K�p�Q1,ekL����k���I��-�4�[{���Mk�����'~m�x���RQ��(ګd��%<�A�~��|E�Z�����%�O�L�N�����Y),�J��S1Y�C+[�S�|��������2���NyBe����5ϛ�� (S�s s�|��i�(hE�A#�#Sv֚z�Z������M�%���M�*�|,�ytL��j�0��������q����哋-B��@_�"M�u�Gޓ�i�=�F��{�_���2��9fM�W��BgG�x;%��Lz�6f�C[Ra�=MV}�k�<���QH?R�{`ɖ��e&�� �r!��M�%Ѐ��A��%~�@�7]ݻS����Rs)3�ٽ������3���B<�;��S���bYvfɠ��o�����@bx�Ұt��ҔAR#���T0*n�s��[V�q���� �:� �h����}������� �[EoQXV�g��w�)�MN�#�FX>��,��h	_��R�t���k�*jw�����
-�º^�6La��Vl�����U��k���r$�P��i��4�}[o�H���f�t��"�G�������(�eΜ!���3O�@�w·B�m%�om���ΏU�㱛����} 3�|�!:l��tC�ʊp�i2P�ķ!�ypl�k
������Aw_i�EDrv�c���>p�o��*�	�	%BT�8Hw��;��z���S����M��I�.�D��fi�)�9�CZ�\�5���z8W��!�%�Eٿ�_�1eHi��/��\J�I��,��q��d�Æ���5�U1'(n��k��� ��ς�(<��ׄ��Z	
`ã����Լ)Tڌ��?֐�n�3�ݱ�ST��G��?J�?;v�F'H�;D�8��l��2�C�*�)�&�t
r�l|S��!M�]�FAn���la�qW�yS�:�A�
6�geOEG�h��*��P����:���Akπ�_ZU�1�7���8U�:C��^g3�N�{�
Bj�OXt�P�5��ӌ����0
�w����^C
WI�8@�P��"�h�~�~�}p5�cB������'�dX}e�p��-H���_jؖR���#�Y3��d��uf�E��?��Ѡ���/^D�@:t~�72���釖i9���N��!�n�!7g~�/��O��Ǹc�,x��/�2K?��U������!���S�Z�&~:�^��(5�<���>��z9C}�)�	bq�̑�lb�6��h�Y,��0c�k��-�
d�N��&2�O%3�[c�����l�N�1�e!g��E/��h���$]����v��_TH�AT��EA��M+�L>�U��NxVS�1�P�Ѱto����d���׋��0DU�|�]!0���d��W,QoԔ�EL�oF��M�v�LnT��I)ڣ��L�V�d��W�S(v�Q��LrM�^�Zw2��Et�j�=�k�X^s�q��`��c�w����H�o3���v����R��ǌ�*֝��mpL �Q'���i�n�*KJ>E>}"�qE��� �����\��-�Q��Yv���G�5N_�y�Έd��;:u	��b��]�����N��]�!|����&���ڧ"n|�nA$����(���o�hlaD$��'36�69 �^1Cc`���"�efKl�1B�_�
tv(�)��*Z��^K����u9����D��F?�&�hD����R��[&�+%��7R�D�N��&Lb��a7%�G?����^n/��)�G<UC�ֆ<�~�J�s
~p�t���&-L�;8��o<#Sg��٦p�ˁ�^8��G3Q��ư�r��S�ev��_uw��^F=��W"����Km�A�����O��#G�DB. $˵��`\���F��	,bi��`���+�O&彟���^�`�̨J�T=	�l��o����~J@Ҏ)3'*�P�����7B0���U]���q2Y�@�u��Gxh�UG8`�>Oo;,�q_��v�
'2��t�����mbb�0�g���F�KҔK�@Q�S�c.9[��:��:B��z��9��	��+��q�Ho�;7��X��IՀ~g�Kk�?�b�Ԭ32_1����O�=�o�{- ��>wп�wk�2�ȚX��l���|F�Y�A�QAEP�ڂ�9�XnRt#����9�eT�HJ�y�@�F���Q������bv���Ċ�ʳ������%@�5���\5�+i���6�$��W��v�S=!c�)`�f;yaw�%\�\C��_W9����|�jh#ᮟ# ������E���G��D��<̔���h:U]k��a�Ct��K�bg΍����A�&�|c�ŏ�T��g.M;Q�BO��|B��3R�̧��eլ�4)7��`�Si���O��q2���19�@u֦��tL�A
�0�vʺK��}Y¯:���3jh!�G�V���>
Z�e�#I7���]W�)ń~Fc!E�t�.2�s��;f}��"߈!W0}�,xՌ�g��B'�ogp�$�P������4�G=��H���q��3&��l�O	o��z/G)]�@jz�1=,�8��H��<1@�����hݩ)���C�6�1}>���<��BZ��%��	{�~�Kq�ƹ|,�hm��'�!akc
,���$�b�$e�����/v<��.��XE�Q�]����q�*8����m�^j��@0>��k�ƣ	9I:�%�k��Kd;I>E���r�%c,�]KaT%�L�;�O��9�2�^�,�@Ł?#A���;��yC��0e�f�O��yfkV��'m�����'��2�{kQ����{��J��O��e��lt�r0ʶ���j�����DK�aa��+�|@V���eW�QO,��ݿ�g�;b��q��&����� iΜ�"�P.�{�_�1�7�m政G8$�g��3%L��>
���0|!A�ȡq�	I|���3�th_Ḇj��{�Pa��y�Aj�.���l���HE�[�ʷL� i����:��	�2Yp��m�$��ph��c94����p�8T�f�� a�U��~�$v��&jӑpH2*ZrB��/"K�k�_�a��H�-�^���i��X��!�m�=4�q�?��3�WsYB���d-O����{���1NF+p����{dVJ��BC��r�t+��Ď�	k��]z��m��h�������t�D�"/|��&��H}�s�j�͜�6\౶��LQ�1�\'RK�F�`+��&�r���hg��vzk��l��!��S|�B��y�R�&�L��iK�yޟ�I�`F����eXWNT������*׽�5�	l	5D3m��
��:V���/�W��bϠ/����s��H����J^M��dV��X(��|��2qI�C��Rauc������OeA�L���Ӳ�ҜV5�#ez��"�ːEE(f�S-�8.��K���a�y�sص@9H���i.uѼ���*v5C[����e��\o��4�G�ه� � �qq��|ㆫ�p"O�]��e�ͤ��:�{�C �sGg�M����M61�N�8$I�؎�=p�7�}�p�� -�@������ZC�r����[���(��(BO5�B��S��"5���7S��l�6���+f��Bm�H(�i20�QO)�@� ���L/�K؟��M.֭�,����uy���ިh9lg�w5�$�&��h_�؆g�b̵ԃ}�{A:�YMA����JQM�ی�~[�/�=K��3��?%ϳ��8� D���L��Wk�.)�_1>��z�mx�}�e���.��A>�'� ������d���Yp�"j�?o�p��܏Z�)���s�$I���	�d�K\�*��j!�s�� �[ĝ�Z[bk�����Va�Ԕ�Dh�.4~����YK���3��~���<��kn��kY��q�jƧ`�+(���[�{��Hܱ���g}��%Ⓐ��\��i��.�}zGZtzk��}����IHޯ1�B?��L1�ћq.�2^�^�!�dyt7��篘��K���P��&���?�#��^�\��pwF�΃�C7ݒ�|��� ��Ne{��NƂ�bTx:��6 ���9�J�h�l(�R-��m=��"��g+� �Z`=a���s���0�� ��a�m\L̤�@�;-�n�h�'���X���Յ��R���4�d�$���������[7�J�X�~�D����JU}�W�0���Y}v'׈�ՠDǉ�A�
��j����|�)1��^Ln���j���HU�F���!E+ɱ���x~�F��� ߒ��Pbl"��Dж�c-����V�X��݈ւЫ^�U$�ܭ��C�����n-$nnmf�ʕ�a��0]L>˱ZC�L@��z� +��g\7��1�)M'��p'c�7Y��ۘ�˹ 	"B�Z�ڧq�+rƫ�L�N3���J"�G�~�Z���Q�|�A�{�}�j-�%�r�s���ã\e6�����!�T�ex"�<�-l�&�*:���w�մ8�9�K>�ѵ��G����ceT�uo���ZűE��»-�Ο��j��m�����r��Os��	��%�� �20+��b�7=	�\Ps��}Y�6��!�3[���x�uP[��^�x���\�����]%}@8ЪK���y bn��U�1t�rWٵ����,w= a{�g������$��@�O�6L��g�>@����c0u�{��� P.��̟�PdC���5i�]�r�KN�2�����toO��y�Ig��
��$�V��a�ܾ�Hx��_I�L����I�er�
L7)��5°�< �Y�W������ڌ�6qO�����nN�� rIrV��0�=��Е�~�\��`m?h)k10b�����4_f1��4'�~'0.�$n����]�5�qL�0oh�y���,����{�QN^��,󁕾\�B�����ϓ�oݸ�Z�pB�����=��>ҫ�Oms��;0��+�fP �W���q�J��|L����d�t�B�f���H�����G��%A�����K}ш2Я_F�������E�ӱ+<��n#���7U��TP'
DRIFy���_d%]���vM�P�M3lK�UIUhK<�����R^L(�����m�?��d&1����ӍtX�$�U�!ф��+��da�'����P&h�?�D����y�*�'4�������ԙ�`r�p�au��@By�jK��B¯F��� aĺ�D5T ��Uڋˎ�>����~�LC�B!�.�}aY����u<�y�������,}��$�W�����n���멊�G�U�6��Y� �k9�|�撀��(K��I�a���.L���!m;�wI"��u�rY3a�*3�i�RY�+�n�A*�7x�A����-W-]�[��f�{���1�Z�Øeg�4L����)�R@J���2Y�Bo��Z�G��X�U���8��=�9�H�c��Cd�=h�^��6�P���9>�TQM� y�}�hX
�s��-�k�/b9� ��$H
������l^WU>�WdNo��S5�3I='҇�bI��UR �fJ���:{8 �����l��#�QT!ߌ��si�W��=]R|���~�,=H
,h�q0rN�f-�H� .�I�	�,��N�$|�!?s��WV0'���pvW�U�dP^Ѷ�ކ��f\���1D��O|S�XD�Y���Sb���R����7EV����6��u��d��<&�	Bk��d+R�Z��TA)&�w�Z%{IdY0������������}�BL����ſX-A�A��F���;�9Yz?U$�3a�XrT;Xᗷ��"CE��tR ZN��rp3��(5�F6Ͻ��	\�����E
�	�޽�<�&�/������d��9cV�(~Sm��|�����ʫ����N�Am�'�օ�5�I���B���X�'�������=��l�x>���9����2N(�g�b�rI�Q��=����µ@�P�>,,7�k�&�����o'k����]�4��+oBN�7\��Ё[ߧ:rK���SXC�2�(��M�H���B|\�zS-��&�X��N��1J����y�1� ɼ�+�H�T����;K�����ۮ�����G4���-�U]�`+��|G*��G�#�U{� VL�v�AU��܏ 1�1&���,Mg�z�)ȃz���*�ҭ�BX�Fe�lȷ�� ��t�h2D�b�8��Qڿ���G�?��8_�2A�	��c#?k�]
�S�j,J_d�/�#�ƺ�#0�J��wfa�]X��)���D���YO8��7�V�~��T�F}k�E͆��@�@�Va�� L��3�sB8p�e�ۈ�`x�'eY��5����PEZ���GV~n�g�҄[X�+�����[�d���vCg����C~�ػ�QB*{��@������~ĂQ%#t�O�:5!�ɚ��UZ)2��B	"]x��J��u[�,��|��� _�v�=p����K�"���$\&V�ע�d7�3�����#��/�ԭ���?Wv2m�ɱԚ�S)�t���ۣ��$�"F�2��,��I���b3�i���}�
2l�!�1�_1`�q�k[�q����+UL;�L�a �T�h���}�@ߑ堠hLCm3�C�V&�3��?z5��.�ŘrE:�����C<���^���;L?Sa�7��5;к�Y�9��E����(�
���4j�TVӱ�=���^;zJ@��VpO0�ռC\��w�k :D��eH__�3E$�N�|[D���Q��0��x�H�{�e���N!�@�.;^��4��M�F
'kE�$^3�5��{��-`�5��+r�w00[�2����E^A���>=Qh�-��N�B���q�2?�[�i��7?��2|3�*9�E�=�d�S��n�l�^�0��Ø�5�ttS�	���sĪb;L��t^�D*�d���j#F��9[t|$�*>���`�]�5�����{IL�v�T(cH��Ï��9$00@S_s�q�����e"Di!�*@W�XZ��+٩f��*пbE(SrlXX������o�han�H��V����ۇ�ç����i^�3y��Xd� �;X?ww`0�v%Y̎���9Y�����$.i����8}LwsV��*/�{�X�J�U��C�%Z�<x��(Ѷ�{9�<a^���S8m�����������yL�E-v�<I�5E�������ɱ.<b��Z�GTթ��� »�pD3>�tP9
G>Î<diJ�2�t������;n���5d�\zU�=��{��j"~xb�`RQ�k9ah�hl&��b.����D�9J�H�Ŏ C��!k�7^��}S�Bf��?XϪ��M=�9.)��`Y�įjY\�Vj��'�F�N@ �?��9ߣE���/5��Kh�ģ��N([�;��v����u�r({2�|�z��n��=���))S��E�?��^.zaGE�4! �� �=�x�@0r�;�?y�W9���\�t��r+���Mk���ʊ�:u^�\ED�Bg��㓁��D4�fA�H}v;���E���nIz����Wf��fׯ�O�&.�qj@��_�ik��6�6�ɓ����	Ÿ:���KkO�<��2Ag�w����L�� �����<ɞ��H�V�����O����4�F���z]�����s����Ip?J1�G��z�v_#�Ȣ�#�H`gS�&�I:x�v�2Q̫�vunۤ.��FȖ��z=��b:>dx��1
ڰ�� ��ω��W��Q����N&;i}�|��s��6Y�&��e�F���q�lq�M.��Y���Rж��@��z����dW���k�f�2���
ͩ�2Pv�0�#,U�~*��$v��7̡\<X�g�^�*����-[/���W��Py�~����U�!7�a�l�i�{s8z���Z>{�R�����F	�!��/�MYl/]��:���L�WftkC���d_��7*�+D<����Ue ,��&`>�&lD��:�/Ggώ�B)����iB����Z�]��9q
eg+��je]��p&���m���t=�N�5�`O2-���|c���Xf�dĀq��		LFK5�ڗ�c�& N���?��mS=/��Q�3�=*8�T|�P��H�Y��+j	�Yf�w��G�G�t����F�!������8��A���Mq72t�*2��ٳ42&q@"���:�������(m/��lN��V0�>�$�z��'�q[����C�m����ґ_s�Ɯ�\�&Uq��kE��j�3���Ў�*no���/7ҹ����0v�>�熻\TX�Q��p�)�w����,H�{gS�A�����Q�շ"�(����oXi?r>|/�Z��rP�����n�w��~��	8��Xey��`��(���?���a5�>Ύ���=Ȳm�u�.c{�P�G��k&ti�f��I���q݁�_�v�kQ�J��u2�V<!=$�62�@��>z��`��w�k�cgų>� $6N8z���fL�oG����%lZ�b0���������,=O�.J��ߨá��;�]\,�m���_�&�S��J����n%A���lJ��m�\��\�!�V//�P��J�Sh�x\a&�/�,��������z?^u�V����ro�Z�L!��%�21� ��幽�#����SSduj���cc��,4��r��#��>�7�h#:]45����DB�M<�$�2!z���.�U�
k�䗂}Da�I�3�Sӛ6SUݥ�>�1�DQ,��)U���Ո��@2���I�����>vwd}��_QJz�P;�8:>ڪ#�ز�ZvG�W��o��LMT[I�S�U�0u�^i%�>]fL�;K`�9�У Y�n��Z���,KXԣ
�a[�pf*��
`U������š�����B�?�.�u���7����~�d�?��c�-p��[�3w�5�j-r�o��l����}��؆�J��~�9� �w��ů��s���9���`�Rj?��g9��g#~�oL
�m,��Q�z�r ��Z0b�OR��=k�-�t��6���׆K�%�}��{�`�[�=�t�㚮oaZ���4?������9Ϲ�%UZ�yr��~��j�XX�r�R��?ֶ́'�J��b��l-vFN
�fiv�s&o������D&��Ak���?�R��o&�࿾ÏQ� �i	8��؆a�䩙���j�:��p�8��B?D L��0!��	�Y㹼]��{���oa81��Al�(�O�굽v��jw$��͐����+�m��6���I�(B�&"�@���k��_R���5��
�OR��R@[�֟�{�)�?4ѩr߫�drݍUE�nt*!]����n��H���Հܔx:r5'1ar
oo? �ת��7�Qg��r�#��o���V�u���R��>2 �;5��_���j�5���E�ZWwŶw��d�&�h�=�O�0F�`,�S;�br;%t�o�[��흜rs����(H�hq���%�ov�\�6����/=��2����[�,�  UB�Ƌ�1do^>(����ӌ=��N��3������F�kpQ�a�5)�����ö�E�s�
��d�F���j�vP�J�Z�ep��_�G��r��D�pm�|���y�@bV����5Q�^���ј����V]T�\ |R��o�ک�<o���m1�~�����i�.�F�k�q�������i��aeR��;��L�4��C1��\��/5�PTi���`'��_�G��@ܬ��,0��a=�42�B�(��������@W[fi��x{�V�pLy�������˵w�����5���}�Gr�4�]�9Ł�b�Q;O������1W��q��J����u�[7�>Aa�T�E?�Kp��1�#�q���W�΋]���t�Ι)��0�Cnz-��?�����Ivp��:��%čk�])=�q���ɂ�/���)'�#�b	?�c��#)y͈��t����%��gSsE���r��Z�?�$d	}�Ø�p}��z�V����׳�A���Q��h#�QŅ���v>(^�\},1�� #8I�������C�K/g��@��G�o2���7k���{��{=&���`��ڠ�,��D��j�\Lh9Q]��F:55w��U��0$����I�ߣ��O�ߘk�MYE�o�Ħt��i�J�1T�1��qDrT��Q�0{���G�NyRa
_2[����]饃���Sٍ�p�b���'�,�����޾]�c)>���?v��݊�T%����+���K鯊N�!M���?-Ω���k��U�Y:sk���E�#�|o�]��)���0E��E�pF���F]Eꙣ3���l9|��di�^�]���t>�[y~��!�P��M \�X{ͷZ��gV��/ޭ��w�_���L��Ѱx��J[8?3��}\�*20O�N �C�eI<�"�b!Ű5&��U�*����[��lp�&�gp`À�����m�?w�Y ��>9�`��'��]~�ݴ_u��.�&o4�M+_&A�
'�0JK��(�����'{���3 ��q7��QN���f�a04����To	�����ŒtO,��C|x�fH߱�O�+5��Vx���/�$�À� ��W~��p�̨5ƢkDx �
�\����H�;t��-�.��\�P^�NQT��AgB�g�-V���Q�M�v�s���1��X���)#���.�s8��G�Sl�m8���������e�ݲ-{D�bܰk�ͣ/A��,��P�� ��Bӛ�F4���b�߭�5����x,`�4FG�'��RrE`���b��4:[E����Zq}K��h�u�����E��e��Ҫ�׮�}0ȍ�5����� J�ܫ�Tx��cM���v��-�aW��]t���Z�~�S9��壭\��"���������je�ޠ����T^�:�_*��8�n�|� \�
g4�2rCET~���>bu��?,��3��^Q��D�*����:N��b�-�f����T:T)��+8�r�B�>^7�L�V���r��ə1�Κ�u}�^^2���������o<Tg1$�#T�n351�/%���{�3���)�A`]`�Z�H�Ễ���&����@�$�	ʓP>���>� �,Al�VS��ٍ�@���1d�N"R�����8d"��ؖ�v�6�waإ���K��-�3 !�̏sZ�P.I~�oI�&�N�־P���s��ۇ�F��0��]?�Q�3�r�KJX�_&J�����bM��kg% ����3�L��>�?v}t&��E��_w����1,��Y�;�w$���*!K\66	Jw����0��6} � mE��ZG�.�i�0��aص�?�3�q��y��Ь5w�7��e�#�`��d�V�����bES�mM�K^Z6k|\ic<˜���>=G*A}sx&5\#���7)�[V��s��:w
���C���b&��A}��#�.�;(%�ȵ(�NM~`�T��,�2Wq=ŇqA�K��g�<�?�D��k�L���θ�-��"m���o�dkE��}J)����s��Uۄ�F.f9
���R��s+�/i�Y×�Ǖx5nޘ�̞򏅺�@^r��@�f( q�߭R��0&ǣ���F8Ó�'�/��TT?G�Ǻ�;X��j�@��X��wJ��;�����m��X�?]A������1�N�n/Rׄf�x�̮�2�=$5��kLƐ�:.��l<��Im�<�x9�]�R�7l�n٤<���u��}Ҋ��*�J��W�K~��Y2���ڍbg��=Df��2Y������e�����.\�D�q����Z~al�Ǵ��pA��'b�z��/&�.�,�����,��j:��p�0ߒ�bl��Җ����gI5ҠHC�V;���-�������σ��$��7����8�q��},�/^&jpdJ�,<u�3ml~KET��cjs؆3b�Dx=)*O�G�5�vs���*ML���\v Gi��X��#9��p��8��!~ �����6��s-��ȯ��l�0��Ƴ�^b�j�Bv���	�����_vfOp�>���r`QDks�	N߼mc�>��,���#ᣢ�<?G���[��pE�0�S(�IE��!'fE�+�_�O���m���Μ��s��3�;���X�����(*ϻ9���D]cs!��x��+�j�9c�U����AD_Ką��ʓ�6�Z�f�G!dv��_z֣XQ��)�~")e]��H�OMK��5'����qG�h���V�fmnk&�6醈P>(��G��l��O�..��x�'a�c���"�X3+>gn�wnr��͋�1����?�7R��#������\�MMs�z 8��T�3\>���*�)�n���Q�O6(�3k;
xh9*"e�q��f��&h��R���Bu�@�M�Ë�P��}'w?�9����zG�����EUWq ���q��k�VNDA<�e�
w!�� 7s��w��ˍ9�����DY�N��c�.�B�O02k�	�]�n�`��R^]ń*T����r�����lSnԦ6Ӳ�9���^�җ"q��29�O�_.�E~$��&��^n*��6����P�I�XJ6�d4F�J��f�&ʀ&@��n�t�0�k�	��p��Ԇ����K|W�
#�uO��ǂ�y+��@y�~���aţ�w?���6���I zȳ'�p���GA�U��L�Q�r���eXY�E0�����V�߼ZE��.b��e	�t�f��V D��x b��#�k&)�Y'�dõ֝�L>b/G�߸%f��/��&4sB:�'I? ����7����|us0�������9�E�a]E�Φv�V�ߟwj����j� ^}|�8�4#i�>���g�9��JS������t��� 3<.���@�a�E�X���w�G��{�j���[w��Bnau�����1��^���ى�,6N
ߐ{
��zV�oY`}�+OpH	�!r6����֟�a,��_���5P"�i�b�w�O~�,�~�_�r�WR�������^k���X��m��(
	&���~d�ja�8.y���1��R�Z�:ld2�J�� �
�2vh�(l��Q1�0{?[^l<��ZK��?f�bc����Γa@»SY��j�=(T9o��:�2��jky����e&T�\����F.R�S�zn������9���0y�q5� �(}��U��	�:Up�e:����9���X�I���EՀN�Y�����RW\�p�o�W��*�����R5c�V*��ob���¨��wTA����'X!y5n��z"�cYn�;�O��U����Ԉ�11�`�:�%�|�b�yd��'�גh?��%�S�~[w�t%���=����m+�#T�/.C36X���>Hp账��r�o`z�7����.mK�0��^J��5��h�ߓ'�'��y2�����c���)w�ݖ}r�_�w�Cq%�b�rP����y�|�v"��wiV��f,%-�U6�tQ@��7q���9R>��he�s��иrBVKp{�lT�bA4�F���ǝ��w��9U�d�z�����T��%�p�
��Ʒ����q�1��I��s/��v���x��:���.$PZ��?� <�e�߻�d�h`l��q�G��]YH3�bq�-��`�л�L�&`��[�_��s�.M�
ރ��[*��_�z��7�?_jV�ٷY.����^h���*�v�����$�� �
ڜ�'���``oKt����39Ob%с�|-[�Q��!�:/�Y�@���w¥H��T��[��z���%����O>�\�2�/idُ�O�vԌ�U������}8jh���F�af�[��� �d�R\�YuIVmXw�qC�R����@���W��yPWP��#	��2�M�&��Q�ѡ���H�޳
���ɋ��׻���!mj����)�[�IQ{TD�s�S%/p��
Ҡ��zQ�vo���7�?;����P��s�fǄ��3萝���}�9g.�B��?�4h�ӣ�0��n��e�4��2�������B�E���7�C����	��K0�"7Ⴞ�/l��k:��!����P�ݽ+D"��I1�:ۆ�k�K�z�T�H@�9�{��y�j2��$P�Z	�Ojn)�]��N�uA�%�D Q>�D�~�VR��"�\�:\QEijsF�\�8�$�~�F2D�>�q1�t��?��Ӕ,N���h��v�����b���b�9��h'd}��}[����npz��R�{�sM}&���C�����ٚ��`��	�l�5��½��k�a2�@0ԝ��PM ��@���R�۹�.J��X���T��:�m6ꡆ��r���ڨPN��E�d��~��Ƣv�Eȗ3�U���<.Q�>U�8��C`�^��N�R>���(��fNU��Ņ�h7�-\5�K�X�@�W~�ڏ�j���\s�y���S �e�i�|��{��Ъ%?�i��@tDLv�,aWbJ�u02�}�RX³�3��0�ÚHH$+'d���U��i%�}:�X_�"�u4L��^�J�yv�4XF'_����nҞ�` ��a9�}�~�j`��$e1:Ҩ�Q0R|iO�\P����b��舖�z�찷�)x4԰�b��^�zf���TM���G7,*��X�V�
v6�qu@� @�.�6��p$�aG�����3�0�p*_7����*c�P�����i��7l���"z~������nK��\F�m%}@͈W��[%H]㌅�����fWb��s��B�Ƽ����"~|0�`�=�:��I&]�^BݭJ1�rnGը�I�����GFT���\x]UIo��R�\j�<?(�=rOO�a��B����x����ɇk��؊��f�l�me�wo��v�n�5[�[����(���gh�;���X�x[�'A�G^hw�w�9"AVG��-Q\X�ߪ���(u�:��۷��<�1�s���;�:Ā�Ԑ/M��S�4M6�u��0��(aK �1��p�N}��C�by�h�Qb�j�j0Y	ft�A�MU�����>�h����C�X���� �g���i��+O����V�T����aGC�S=w��,� �@��jH%+�p����5��6U���d�Ѓ�)"�t �Hz����i��ݢ���$�ۈ����Aվ�;24a����9�ǮIu�ڴ�c�\�1�i�|�U$�,'�,�M�nȤ:���_W��&��e�9� 2a�@v�kr}9`�k�MA>1���#z�n�Qw��YO>�8y�pL
1 �*Z����6 ?�$�Zb���� F���7����k'oY�
��c�A�e�D�=��>�8�-�Vʮd��;�����y���#�|� �\��wE�3`�G�\�pv1nyrB�0
���L��q]�@L�/O���+V�U[;�҄/dM��M�t����y$������Lq��$V֢y������W���`���� ϝ���&7���f�OS�������i��g,]dm.�[�F�M(�\���#��Og'�r,�;d�ً��3�����ej1�K��b3(��*� �=��$-��S�#���g F*H��Z�KiΡ���Ѧ�X���[�+B�ʐ$��Ȉ#����j@��Zsr���
Ȟ�7�ks���y�W��{��)��>m/�i8�v��ZTW��٤]���F�Y�-�M�|D�P}��H/�nzm�:�(�s���[Fޣ�������^i����6V��~U놿M�eH@ 0�ML�}�}s�S���:^+�	l�� �����C���H�@���ֺ��d�o�ǒ(��&�-����S�E,���:pU&f
�V��O9tS4��W5��v��_W��R��*7 ���,���b�y�ח��܍V�7oC6��߫`�I�A��+�)�_7��/�1�9km-9_����U�ɜx�[x��z���o&�&�� �'�|���a	��Ilס3%?� ���1}UiW��(=��2#���-��:�.��c��&E^
, A����>P��V�h����	ߙ��l��fO���S���i�@Dp1~������H�h�h�ס���N��gk:��v�.+��I�d~�����v85�j6�*���;S�XƼo%�O�w=��@H2V��}'o�ѻ~Ն{x��v�ev���'%k[����U��w��Mża�%�7<~��s8g�L�6 )�X���ݴ�U4@7F{�䚮	�5�0��fq��r-40	����q{��}W���`���4��QrG�\Q�'Si8H\�����6+�6�~lV5�Z�/�Ϡ���'h��
W��o��R{����\��J�M��*�R�����]���-�{K���x�A�r��A�+5�j��l�W?e�y<��������i�	�EH��~��Y�6��|�E��%R�;>���]1p@*�:��>�?���y��k{��$�Q|@(F\GtV��XY�O��i���&�B7�W;,��nRAm�ƃ���h��b�Mݼ�$�>���M��3ޏi�(��u�`QUm�h����-6�8R����L�@x�@k�xp4!��1Ϳ�s�3�c��\~���9<���ukň+$��"�g=�#�ڙx:����.����2u�F�-�g�=���t�m��8��gA��ښ�i2֥��և��}-��K�����Q%؟�joɁו��a����R�^]6�L�m�N�����O���&��$�N�$���������c<�t¾5�� U�H"����)5���)W��Y�͐k�F��F!YO�:L
+Ό/[F���t�Z��8��&�%�O�r)H/��_&���~CP�Z��_F��r�N^;,�*Q��Uꆷ�OҘ�^=�\�|�>g��a����þT&�~��*�4���Y 7�z�>Y	�T�4`vK(�l������=����/�wHF)q��(�s�3�KB	�m=��]�	l\ڠ�I$�o�,�N{�C
p� �HBͺG�0�/��A�JT�{"�~q��T�
�
���c�����5�X�,�@��� �>n��P�����N_y����z E��&��f�bF���k7~�#�}�Wg���7w�T�a�;
����-�.T)!������%�j�A�q�D�2�]_��*�1�G����� �ǙJ��Wִ~���0��=9�f�A���E$�,�B]�=�>R��#'O"�z�Q��p5��#P��2���?Rv����[�fq��|�!7�H�Y���!�̙d,�3���D�AXQi�ZH�J�W�[�D�V>҃Rk��F�4�3�L���*�	5�/�� cNG�0rcJM���1u�s��$PW�l ~~]6/��x��n��������������7�
B�๱9{ rO4*C}�ݥ
}�)2�(}9�WAr���+��wE��Jp�ྲྀC�o��X����]޸WPT�]1�1�����F�	?�Ϻ�M`L+D"�W�A�=v�;�˜v�i�75w��b�D��4v	L
om��)�?����$#@)����������*��qi�λ�/��툲~���	��|)�Y�.C�$ʹ2�0yX���� нy�vMr��� Oy��@Jp%z�B,��(��^P���.�l@���v&E�ip/���#���ʽ�I�f���1��6tx�C�͏HI ݄�=���_�6�6w�.���`�����-�_?�vF0���ς?�կ��|Z�jc;Ϗ���X~��$9��G��
rl27��;k��z$#/f�(�{�OΆAw���Y�PYql�����n`��������RK�b#&���H�&�jg�����(�j�	A�p��sm�k%+?�{�"mY�e4+N쐋�9n�)�F�/FBT��3��t�D�K0ҶĎ���#�� �Ҵ�z��v�%���X�:9*Y��V�Q�,*�49�m��b�b�=w�oxBD�C����IbH.�H�} �;ꑐ/�=�K߉�%��}�j�:�Ԍ/r�﫫��c�(N=V�?wV��{w�ldAr[BM?��S�}"�m���� ����1�?|��ׅ�ߠ
U�!'����xq�mk���M;�}����F"��֔��FY3
Y�j��Q�P1�U5����42�bD�������L-;l��)o^e��"74*Ã\D��� �5��{��*a���<���"���\\�GM��_v����*�;�?h3_�5,�����H���.-Eo��	N@'����	Or��,(&�n�h1t���P�S<�t��墈\kl`���l�tFx/�ǝc/,[�{��e�.��k���bd�� =$�,��ڀ��t�����i<�G�hE@��]{���/��L�R���$~�1���%�K$��)��lN���X�﷩`йLm�bon�1�W�hX*�A26i�8��1M�۸��s��Y�3��{����ޯI8��Xb��:�Cl/n�ʷ|����6j�S$�����ɉ����P�o����GG�@.�j^��n+�S)���������i�Nx�3��3H���]���"�ғ��UE��gx�����"1��6�=��P�*4�ݐ������,��e_�lJ��~0�ak�+��Ԉ�83'>�y�ȴ�2��<�� ��F bO(@�ז>�z*�vs>���D5�RZb�q��1 )��L����9:���˖j�ֿC�
��Y�������J�����z�s�ÚpZ���}w�V�h����ͅKM��}-��g���P+>>�:r���_����;����?k樹kU0�R��o��_G��'7p9y�9�q3��pݢ�o��s������CE��Ր�o���f3H&��1�g̄�Kە��jH�h��-T��>e��$R7�W��S˽���D/>�~� ��.�gg��N* kUy��JV���.s��WdF�bHg�3�݇��(�#�%}%��q��M�p�cv@�N�Y�
�"r�T�i��BH&��`28hT熐b��'�x0\͹.c�S矰���G�I�~ߦ�YB�d�I���I3����9��ӳ�Km�ŏ�s���=�:c�q���2�y��� D���k��������qҦ��;�&f��27�dU�7#�L�����m�o�(S� t��� Hdk��@O�Xx>��|�шl;-�����8.��B� 9�;��F�A�}燎�������1��q��C�!�o��į�(*�´)Vo?��5��g��/�Ǧ�;�?���9`�sV(���@�����X�HI���$������B�+?Xv��VYo�t�n�n��#��� �(x1!�����V�3L��O�����dF��f�S�|��m&��G��13�A��G�	�+��Fءf�^�6���4�e�)�������dø}�l�o�%��T��W\r�;��ʌ�լd����j��Eۘ����E'_F^}jl�9/�&�Z�j��ހ��j�i�f���=_r���ߚIl_�?t�؋��Z�mZ�>E�Y�N��Q�#�/N��]8ں�zR3�\�r�Z��)BV�@�o��ٽ��QE����#b�@S�vEU�q#��P
�����������'z�#��{���"��F_�v`�8��d�[h}I;�U��@��B#>�Lt�P�e�W:��~X���,��R�.����ͫy�x�>�T���������'R9T��ˤ����,�*qo��� .���h؍Fs��"��eX��o~W��G�چ'�և^����	6e _PdN�j�R����0c5R���e��<5j��)�O,�����a["闿�ui��K�T��J�˔����U����0�xW�<!R�6̝�@͟��"�G��'03�����?R�/����!8�i��"�������n�#>{������B#�ެ��明пi��v�����Zg[���]��֡7vm�9Ȋ�5���������d6��j���Q������d*:$:���;��|)K�􃮥�z0��Dեhn(���L�QS�o$�"W�Ԝ�Ė�@�};f\�6�#YK�ٰ&��Z-�}��I�ź�ͬ���r�p]��tW��vSy�&se�gR�S���I/�t�ޯ?�������dA��u�TJ %;S��`]^��s���V%fmRp� B� x����5�$��lcv�6l�Y��D�*5j:c�)Cg����ݚ��yV^�j�#bG`���������+K�hn�r��./3Nl��%'/9�"��.�WI3�L��C�r��d�_j3i��3���P�n��}�#f�]�lExZ��ҡK�M��2Љ�.�j;�Y��nćME�_l5�?(ԏ� �GI� ��F����@	�<+Q�q6�D6;��W�2x��J8/ě��# �4����K;��g�ٛ������
�6����0¤��+亅�F�L~N��os���r�i3i��+�0{�f~��I��7�b�H]4n*���SL�(
'
a�-�������K��%��|� ����v�^��K��Y�a�u=[B�^�t����k� ���̟$0��ˋĴ�xF�i�W�k��0�egKE5E�����.�W��֦v�mk��ܱ�aA6�*�_|AK �T�C��~�'�M�珱'�3�r��6��t3��B�w�������X�H��/t���4�W��K��������Ѫ�����M ������K�t��C*}sm6{�����`���X�\P1�%"� /�yo4��Ҡ�m�=m�����xw��)=�c�?S�	= ��s��NrL$����`�7 �E:��ا�#�bbqylYQ�7ϳ�A�v�|I��2ˣ'��rrB��_�4�qa"�L� R�/~��HW�Ԉ�B��������}��w�~}f,�Lt=�>�jq�����ˣ��(�\�(3>���NuC��+;)��y���b�W�K!A���za�;$EK�����8���Yм̑nɩϖw�*�����pj,8w�F������ݓ���N�E`EJ�� +�����A�0Q�
t��t���C�5\l6���YeÖ��V�:���v�S��nP8mm���=u�,ìF0�cλQ!��|.�1�~�8���q��y�i�a,����}��ē	TT�=7֣�PiݍM
e+����\�	{n�;���Z��~�5�+E}j+Ǝ  zUs��aS���^���x�����u�x��%0 k�6�������؀��=�R(��a!�$BVU���	B�����Xm���d1�Հ֓�B�Q)(a������k���3#���r*f�V��Z���f��?+p�X�$��ﱽ055�k�%�M�K�G��3GH';�O�P�����n�AkA�1L'X$�v���\��w�a�K�����&�'�;���9���O�<N���I��֞s��2���V�\�>�
ٕ����;��ed�Ԡ�4�o�BBfL.99Ӓ���;�R򶸔�J�#I�=u4�+�)6G�/��.	�L�3u1��7lRվw)�g�uZ�zS �F
��9��a�����1
7�l8�~��Iz�/0#g���W���6�A`�5Od�!�ћ�m��B���kS�����J�6A�1�ŏ��P+�&��֌��X���Qsɸ����@I��#7=����^�x�)�\�v�Q�cj5s�p�	��&�����AP�v
r�p��˨_� ��ٌx��\��܋��>�d��`�Р؀�K������t�j�!d7�.K��@eO�f����z�J�����Bt�$9y����Q�4�f���׀0 >�LeD,9<�nd�� *lSٽ��8��1�M�|�\����)AS�ju=�G5��}߇��yW�y%�d�
��6΀�Q!�ͧ�I��^�ˁ]e���D]�D�.- ���oݮ�4?Vج7gW�����"yqZ�-6��<5�+�q�'TabDCS�d{�\t�Jy ������m��aM|b�w�IN�U ��&�h�pn��;²��$~j�,�G�/�)U���k�>C�NDӊ8���Pa'��ܺ�Řs�b�cL0��\�d(�����❖�*H��
BHO<�us>;�挱���a�v�ˆ2;k�u�ۯ�yd \���U}d�m�Ic�IF(�R���c��ƌk�Ә�+�6D����30�c }�VU��>$�g~�.O<\�u�
-��KYg��+!y��Y��wV����2U_�c��-��nm�|��+Q`�bvݘv���:��Rl���*o8�^��<���ڒ0ǜp�Ûj]�{��>�q׺}��F���]���ǳ�Cُ:NVY���l����ԯ��g�Mx7GBQv��Ę{�ctg]�ȍ�QIV_?�t䉔���m�J'�봡��!���W�#<3ʠt����]Y
f�P�ޏ��\��0;V|�`�Aa���?��}cDϭt����"�&�%W�0�
3��4ݩ�e�V�T�������*N7�|榭��:�N.��h��8���_�ꁔuܡ��78L������D$d�h#�ݞ��A���v����Y
��K�:�x�f��Ds��85X�:��j��b�P5��r*���'RUI�����"b���j����i���z��m�toR8nrGn�.<�#��ٛ����'i�<�#>\�)!���}`�˶�[TǍΘ�E<(&�,�.��@x�*���,b�5�������;�BZ��C� *��(U^%�n�zs��P~	e�>��c7���nrw��zE�9�P�c�I��#׎W.$j)�)�������c�8��z�Ͽ"[����w��1�f�/[6�\��tx��ȇ�j���ģ2J�Xr��iAh��}�!gYګ�����*a�D�<
�����Q�ds�6�Oء8h�q�f�\@����	�8c>x��%[}�2Kf�M!�xy�L�^����X=�6D��r�XR�7����-����	|��<Q�GQ+[��5]\یt��U�9|c������HB�>�YT��K�z��n� e0���G7�ln�����t�@rC��J��L��� ���GGjhg����k�,��v�����<�?M$�����z��EM&��٠6�Z��a�����!*�=�8P%_�4����������	"����'2��
_%#���t+*jĕs�,�%��ƺ>�"s�s� ���"H����t�K"Z�0j�R0�7ۈuJxi�X;�"a�s������Y�V��LS��bAW�^���2�R$�#]�j��Kϕ�/3�9��c%�ƒݕ�mf=�<����*��&�c��e��:Ε\x��!$�q9W��ྒྷ�V_�8/q�3ls��7�+XQ�@T㹑��)���<��ԝ鬫wLW|��l9+�~g�A�'NS�˻QSk(��X�@���I����B���'���{��£�Z�jM��I{���*����45ha�A��r��:'G���YH�^�3���D����>�!6p	��G�_\j�L�1Cc���E0�S����x�"���(�W��r� b~ �p�Mj�K`&����=tj	�9��n�sF��S�{f�#F�ey(�co+6o��C/��]��O����qQqm�"�؄����7�o���4��]O+V�{��Y��$*6��rC��6� �~:��rM��G�{�T��Vu�86�2`:5?u��U�ѥF��k9�d[m���9�7'/Ԍi��W��7��\���_&N�����(l���oi�P���0_m�����T�W���k�~Ŀ���[��EuOUr��1n<g���{�y�����_� Xi�!�'�4԰�_��'DK0]��H�s���Lz:Iyn/u7( 	�Ew��&�r��͉e���d ?D����?�%G��GL|���ܭ��l!���Hw������Yn���o ?���b����2*)��@Z��-��`̠����#F�u:{?����U�<#q�uF�^*�q��O�GrZ3;�`���|�����۰o��R���:��`I�p&���&�2��g�������2�Y���1�>)��OsǙހ�'�W٘�tY$f�2�/°ڛQ:Q�6GNʑ�x��v� ��&\O�C�$z���{"/ːߡ�Ɍޅ�\�q<���@q��}��裵�!n�� ��v�}
��<�?���:���R�G�w�ݮ�1�r=	d��Muk�z�l;�*��B���/P̌�6�S�M* �6��{]�����A���1�����o�4+��~
�N吏���^:�OElY['b��c+i
��
t#��̪l�c�j��rF�yg�.ϧ)��i��O��v]�ҥ�����)3sZ�J���'�c����W��G��i^�RH����u��_�Om節��9�Sk�(I������Et�*���%�g{�f�­NR*fp�v������U5}�9�=�
�3"�wn-����v���p�!R�<?CXӈ{�,�H
��4��#7QAi�&;e=�.OKj&������!��T?0=�O�R���=0���d��4���i4U����!�8<ݸ�����[���X�YC]\�g�����q�Y'F�(^4�$Cq��p�r��^�a��~����@sZJQ�QW��G�ۉ��W=�4�vW���I�@�pr���+P���r6��GX:L����^%cp�/��!}���I�mJq���pk�����@��P��?~�â�q�,V�Na��w���ͥ~O�W�^�뤞G����N}~MJ����]Tg����ȼ,���j�9(����mZ']��s��I�#%r�C�������f�H��=z��9��@�B`:���%
B��,�ir�_�Y�}���$D��z*_�-dY)�2�fL+{q�{6H�0�s������(��`'}2`�
^���� d�g�����;��}��9 G�BYu .�b���jt��pL��~�N*�J㹭�#�4l%:��~b�%�/fE�x�R��GO"�8��=�Xv�~���VK��a6��/�?�o��$�7������b�U��3J].A���(R�K����;yPf2�s�0���{����7����#�_���n�'�\�d�ot���S��/6Ϗ����H�U�4w�	w���G�y���7�t�����vv���5zkym��t������B��)~m$n g�*h0�k��=��oإ.�l�z�����-���x�� =�I�L�K��Py�fF���yB�#HR�|�l-�?�4�t*]�@by����5�[C<r>}�"�X�ϐ �*|�Ԅ�J���-�~ʸ|#Pe'ڮ��|(ϳO(�x�w�S�%�ռ,��1e����#<�I�\�����Fǲ���B�9o�kc�����4�i�k��V=�NnLv:El[��OC�x��u�a��a��>:9mL��~j�j��E����2�>
���u�z'nI�*摾yj���Yh�s����Q{݁�as��X�-�7*Ph0�l�{�s���f�nV�j�)�_6s��MR-ʏ{X,���Pn�?������bW�隽�0����ؠ ���e�{jB#0���U�r��:[k�	/�s��s4b-{W��Zܨ4oA�@����Tddw@�~2n��o�a��<ښ�Iu��/3g��Rx�������He���Mϖ�!�� ��x$ �O֘�b�j�J�ˊ���O�ĢG�����6V+��u=��j`bb���*����m�P�؛��y`l��*ϩ%7p���E��J��X2��z�2���R�C��?%�f����v\�?*�Эau
P����<����J����V�2�ur�Sa�2��o���:���!x�H5����4��R$z�S�Qٯ۠�$�H|O����V���
���n��Յ_`O�|��
��g4
}F	��F�����h�}���6�dF/����T��,Gy�|2g{k����;DZF�ǔ�j.ދF�`��Pė^ԍ%ͅ�`r�w���C��	���&�fo�`�Ոr�,��'�K*�e(C��}.��=ƻ�.'r�SK#9�!�y;�A��?�?���<?�� �ɳ�!�K_?�bB:]�i-�:���۷���p�l7�Y�xB��摣�Ȇ+Uq?��o��_�	,D��[��J�j�����[?��	�����ʤ���1'0�7!\^ѹ��| :v����V�\�KVY(�zh�����BϕT¼#��J��ީ��M����)�2�6�%ٿ�f
C���AmwJ%�_1��X�X��A8�t��y��o��n�4��AX{�]�CTަN�,7����<@b<��C�"Ċ�'ȩ��Jc9��E�u
�l�.a**.�\Vλ)��m[�|��j�{��7��#��|x�ăǊ�6P�$�lv.yj���SB�������n�o�wT�]4�G�Xl��<G�! �#��������M2y1��6��i�W�,l���<���W���,2d7ҷ��Z�Q/���d�EK�� �����A�@*ԛU2e�bRMa�=?�6H!���Y�7���c�����P�����e�T'����@.F�L��O�'��?�*����<���h��W�a�4���?�bz�Գ���4������fɣ��_��t8�F���b3`K}x���R�:QE;6vT����6�O�R�Xc*��FT�ïT�Y�g¥l~w_�Y�!*:�޹|���WX$�u���R��LX">t�۬q`�K�Zn;��l�9�{Z�'����彊����ჳ�ʦ��Α�( °g���.D.L,ws+0�`������(x"�|��`B:�62G�2ۅj�J2�(�f�K������"���|���Q\C ��|���aX]5�,��Ļ(mő�gn9�!m��X�Vs�L����j�+-���O뚘J{��{�!����L���:����- T|��7�	ϫ]��T���U�zN�//����<Ha���|�l���e�=I�_�1�~6�D�q�'��{�/�#� ^���a#,�{x�=n�G%���h�kԡ�����/�m9�ԟ���\��+J�	HA�O�܁��t�%&�Q�!�hq��S�8�>8ípҌ
���r��v�G%�c
�y�Q�]�$a,�sfr�k/Z;��8Թ��;��R�T���}��N>�|���Ԡ�0Ij�������`B��!�=B���A�Z��O��ɚM���k��� �!C�;t<�T�ױԋ�$��r��	7�����Rl��J,,������e����4�H��BZB��Oh����4�ZR;EF�z��	�J�0?q�����ʐ�1�����x]��#�;�~.s��e�Z8������ďl���������!�w�Z����D�/�8F��S���5�$��P[�1�΀��g��v���:uI e��k��_���+q����l�
�bM��)k!���s��0xv%^�N��H��k�n���
����"lR)C�%�V��}Dou���b��)�].��8Dą	��� Ѝ��n�oc����j}|�2ߵa= �x@�F^�R��|E�`!�p����g�sQ[�Q�q+�C��׎#�X��,$_�Э�
��\�uO���o���Td�[w���P�!���S�W�	ݛ���S��3J���� N���|v��cހ�ٞ��z8V,���[2O��ݼ�<�>���kW涒��~���7�e8��%��Jeq���ÿ56h޸����\�2غ�`vkdðP��N�}Nkq���5�I�E�F�Qܰg{V(������Q�t.��!�м�=P;߂�kbi��*}�$�r�ۣ���C�6��k��h�!!;C�#����nl���`��L����U���#�L����j���m[}�(���t���)�����z��g�P��)^|ܥo�� ��iL��M7rbhXk�^��9�w�w�8�~�0����uJ
P&%��X���p_��n1.k/�A�f�?v^�˖��t`̝}?plŁ���2^x�:2)���!9�c��|��V��o7=��xả��x0.�H���rO1>^�'{�J���1?\�ƛ�3s:�^0�27ќ+�8�5����gب~�s��������/ナ��裦�͸)���%�P�I���>f	��d�U2v�R�D�T��a�i���}���=�e޳��#h0��d�����􊋒��s9�B���,h$�4�v.(:�H%�Q�L���"~��P|/>K�vk�x�kC\hr��٣��#.hi�}���6ۛ��
������p��нսM/X�EȈK�s�!#05=�1dX}ݮ6;$%�I�x��,�We�ɿ!���PK��l�$�O?<vJ�4Ŏ��Tq���x��+%H�2�ɳ�m�"øC� �l2OQ#q���zn{���=��V������-Ƨ��f`}���[	��VY΁n��*�R�Xt0Of��.�2�9�}}�W,���l�)��C �\�R�W���A�z��3���hm���m����׉Yʒ�������hr��
K���#��x�vcD_�ܵH vK!�5=J=��#�4sh��>�d7�6�\�����|H��6��B��Zx��'�5ǋȟ�{�r�L=�sw���zzL-{%�ƹ�5@����hx븊񤥳N�B3�߫��8�1�g�T�=��P��h�kx_������/��*ce��5���j�De��fd3����y�����z�h5��9b��t�T�����4���AD����T�o�C��y,���2i{�Ǖ	��Q��ݘ	�c>�87r% <8��эdDpҔ�P���%zӊ�i�_v��SB���wiID�2xE#��U�Q��A��`�v�<���7�+��Vu<�x��=�Gުf�̢�r�n���5wᷨ~rhS [��
Έ�_��@��3�g�����tK�6����P��A:BI�|��ɤ�A��]?�<�
�_O�{�C@�M�J���㼊�+�M��ґ0Tt�в޶;�c��_ļ�������>m�n��K���3��E���03Zc�z�Ԩ�W���)�2�:{"k�pU&��p�B�������U�@��ʜ�v��3Ѣ��:R_"�˔�t��K��(�y�����n�]P6-s0� j'.�P��w��b���&�>���dcl�BNÜ���3pP�`Q�U�;������r�t��=w����ٵ�0G�'i��d���6�$R�RI�T���)Mv�Z�QޙݜA��S1,�����U��fy��#�ۃ��k΅�a.���N��F�12B�&"�E.��C�-�Ȱ���p�׶�S�tn��T�q���YTA�SQ;���B{�!1ZՅD�����:坒{)�s����I
1X� ޳$6�����g��Ζ�B���
F�_�)s>G��2J|�������\G�������S}x5o��=<�5�A�n�����r�0�}�O�θ����:z�YM�����;��75o1<����ס�$���K'<���\?Չr�莮��������5La&�B�������U�',(H��;����/�<��:�/�䪼ע��]L�c�k���H��G����Jv2 �i�<7�D>�;�����o�c����hS����k��Cx��?9l�j��tpW��7���QL�ᆆ��_os�45�d��WF��4~�o�]Zru�}��o1܄���䌈�HA�!��\�����2ȬLp���?�B�n���	1<W�~I�S7�9����;��+&߁
��f�W)Z~�{��?�pG�	��Z�<��N�@�
�*  ښRRz��P2��צ��DDp��VX��*��ó�������*#�O!��o�'�M���*b��]�����"16O{�iUٗF�y}�.�B;��������:~D��~q�.���9�ú�$>)��������ə_��;7V�O�~�ke '�"�w�8�<Q�RD��+��c�<�m\&� C�U�,p���i����T��2.f[�0��aus�;r�-j��l�UI��r�p<��`n��7�j8�6��Xs��i��h"��_�ĿbٽEȡG��7n��w�xf�������X?���D�
u��Ǹ����>��\}�A���.���L�i���=�1�/|�^�R�B��̸�����f$�T�J���qp �DG�X����4��g�X����!�bl�$7*W������]L"K��VT��m��-���P�/��$�`�ԙ�^�����5{^�0*�y{Q��N���#�c�Y�� ��ώ�G1�;E���h�/p��;�IF����^�6�Q��׺ �̙���a���V�SGk�" -J@5����CO;V'�J� �E���M��<!0��,H
��|ʬ�PhYv�K
��+0�]�+Ջ\-ÃU�gh���a:�]𲍙�.$�s�?d9�}'��ɩ�Ƈ��
��F��.���e�����"N�W-�[4�Ϟ��r6��Imb��Jiݲ�q9`���B��������]���$Z�X��&�J� 
���r�ʭ�H�_�Op��l>����{��:���
��N3�a�<�m���~����Z:���\��~L�uڷ�@�"�F6��!L�ҼsT�����4o R�3z;�z��P9'�G���~�=&,�	*E3�9�4k:T���>3���۶��f�����*|���]7�BC�����a,|l?�ރh��U�A�3�oھG�%z�<-z��N����l�|H^Jch����g�hk�'�$����>�ֹ.S+��-�#31�7i��^ݖ�'�ԟ�jD�Ĥ���|_�ϽiY��bq�{ۭ(��P�Y?3rU��V�+�+=s2�Z��M��y|= :���;Wl�B�}�S��r�ت���?�<�l
�Ww��y׉S%�Q� yۦKQ�RB�<��o�h�%�Zfȷ$�m)��;~;�/:�G27i����ڬ)�K�g�rC�&{N0��Z�4�-$�K��R��T$��a�� H��VU6�.
kyT��:�@�T��]��]d�}�R!�J�?�Xc,<+��FJ�^�'�5_I8�?��Kx�e�n�}F���F�Qތ�mc�9�rC\S��t
��U�B��u�����6<�Av�G����
����T�<C9}�Kt7�	��t�9��F�yo�J�������od�p!�#L��g.�v��͚���^|�6��z��e�����K4�6U�c��`u-�[�xlW�VܤQ����/􆗸��n�ڈr�Vdm�YLؙλ_&����@�l���0g��PP]�⊗�	%� bB��C��"�k�E�iI�3^2%�웯G��lT!�����U�F�����p4��
�q����y`g4����H2���	�����7�K�b�}C�Y�/[�F�����l�m���N,���x�y�!��Ցg������r� %t7y+Ļ�zM�X����S ��0ހv�2���tn��)/��P� ���ؠ�-�#�/Y���^�i{�!��x�6�-�h
�M֘v^w�K��WTΚmu�j4��������m@�TayI��Y_w5�B�:��G�DYz�Cz�ih��Z6��!��ii<]�ryC*�4X�Sz���q�:ԦJ�UO�����E�5��7I]��F'%U\
�7P/�p
#B;B!;��JHZyX�V��>�r�N��d��ж@�G�[
���XΒtu�䏀sx2�zJ��bi�J,�S�\�"U� ����)ԖU��{����\���**n&Z7UE�K�f�T5��[#��l�I��X��f]� 4�M��̳
o�ҝ���k��)	Om����T�RA�ց�Ė6`աɃ�Nvp0$�Wz[�t[�"�@�US�I�d�6Eg��i��>�E�������ļ�J+�ܖ�C��b�ߊ�F���`�[��׹�m|o��.~h�s�|%�*s#�֞�#N��a�*��]`,�ΦD����P�ŝ�U8�Y��M��<'�l���{y5� 1j�e�?�f^��&�~TU0`)���Bj��x���F|�QQ�^��=N96�o�<�w�}R�Ik.��'�9�o~lq�̦��
Lm�϶*>�8��َ��{q��E�"���� �}��}����<�����]��V�\�aB�����8�8�����F��6QZ϶su1,���m��#� >BQ�.�����8۔ѹD^ٴ�2[�:$e�&��\pS�;����}��V�)U����/@?/lE}C����B��U^"��#6H�R�L�?��^�}�j�=a�-g�otm/�yQ�H����������h���O��Gx�(UwU>e��D�"+��j2[g�ΐc�C�����F�(8�ii�zr�k<��[(�#�6��%���~�,'�QX���%��K׀�w��]<�t�I�>�����ӻmA�X6XV���療;A��c��86����w��!�^?4�4|�h=%�-bX�Q(
����e�2c�Y�y����/߹:®��	��Y���#�ڻ%�ŭ�f�eXΌA�q[�#P�[I�K��\�-�늗��*xX��~fs�a�ܻ�o��{v�x�v�l�We�Hy��sI$R�zj߃X˅�Jk�s�o�a&�+�N΄\�K�e؝'nEeY��>���
]���h��d9:���7�L���D�o}�~�pv�5h\���-�
���:��ާ�?A�n=��q.� c^���S�?����~�i��췿����9:>5�p�C�lW�T���o�%ȍ�F��[)lt��w�`�L�U�B�G[���ㄅ5%VS���rp!C����1��Y�xD�z��x��w�P c�31&�ǃy�&��,xL�1ȥ�&�(X�#�{ �p �]��j��R��U�)b�5p�)�k����@�a�eú1��`E��mt�&g�k��s�Kq��{���U���+Q_��F.ZoА��w�\fSL:+&f��G%�Ԫ}�J,�VL�^{ D~���VY½���Ԯ�4<,R�*���jB#�q����+�ʝGD�NC��0�\���_�-�3����S$]R���E���Z�T{r����z��~M��GF��k���ǒAS�F��l{=`�*�'3�����j�ڛj�n]���5�8oáQ/���%�$/Z�A兲��GZDͷ�!K����(�Ӏ��K��s�4� &�+�k�X�j�i�=N?�z��R��oƟ}Z������VY(���X��h�E��Sk)�����'0!�Ġ�Z�����������޳���%נڈ�;���(�?�!�y)��N��z��H�iJ�״c<��~������0؀���슆}n�r��`q�~�V�+�A/���/�k>�^�o�m8D�����/U�&��]o�G�˒��(�\��y��6H7��?�[���(��O�.ƹɗH�����F�Zo�d��^�?���f����\l��Ǹ��eA�{���dj��D6���c��*)?�1���xQx�F��� 6��S-�<vVPd������¨�Ip Ěý�+d�M�R�̫����g7�#vD�1ʛ��mкɁ[3�Fx�{�f[�k!5�T�V5�y>�n�br���l�pX�)�������0���3�Ax��ɚ!�q/�����b54��	9|�'��?����lbҊR�:�q(���X_da)�"�R<�����Y�,��?h��w>Lo$B�~s.N���	�	�F�@��p?0�-Ku!��(�u��u�(	]�e��o���jS�h;m�K�Ht]���p���A�����1^�R&�E��q��;Z�����Zd�튨��ZJ��"����ݩl�e�Y��2�90~�� ��Ѝ_�>�~���`�K]O��F����B��j�ĐP�4���{��'��[�s&���� ��S�e+�F�pqi��>q���R�=.N�7�ir�q<c�H��b`�T+r�+$�7�c�����	�1X::��~J���Z�˂�����s�!�%ޥ�J��'Ң�x���8���4
pD���,e,��l����'��=1�sG�`��7�77�����׾?�����ǵ����(��"$�'����e�cCVd�Gw� K<o4�ǉT8�{D���1LC�-<�������0�>c���Ո�E� ��oIi����u6��t�H%�
դ�
�ɐ����J� Ds��O7a[�u����C�\�Xzxgێ������y���qk�5T0/)``��J�ఐ�~���Җ���O�tU��5�ZM	0(��3�UBQGe� � 6#C޽����ͭ����䷛'��	fp�$VB�y7��C�Ҿ�#��Y���D�㉊�_�C�v�AONb���oo0N��]��JcWh���fr�è*< ġVV�LTn�m��6��0���С^{�!z�4F�l%�K�e��{C4?�Z�~�^	���[a�p�������<��b�;J*�8M�Qg/a�����u��11X��]��nx��Aw����'���^���vZm�F�����/�e^���/�M�n�n3Һ���^����L����:�?�##� M=0�.k��7�:��,��T]�����+x>���"�����#��S&f�U��z�4|�e�R|D�P�Jk�Q$	#�i�[*Z�)d�;��*�>zy��S�@#%Q�����d�\a�q��?#ML8���#2WxS�J�u#=8[�[��
|e�܄\G�c��|.R����F:t�٣��8�_�H�3�fc�,��!��>���*d��UQ]�愣z�>*'R��A/�E��l����r��C@�mw-��j�N�:�Vg�#6���4�������-�(1�ZLfT��jD3b�4�Z��L����Ŕ���0++�cvb�SF��b`F�q��c"��%H2f#�tf+c}�5j��Ơǜ�vA�M4	Z	*��u�\oLN5�p
7��+�sC'r5D,���k��E��*��I�B
�1�E��2h�="�H]+�2ǳ�CO�6���F�����ׅT�W_��<��l��Tعlj2>W�$�C�W?�����.�.gn�Ӥ�0�(��cm�ۻK�E�%0J�U���,��C��IIbs�^������/�*!uoj��A:�ѫy
��ջ����rッ�e�O�Z��M4Z9������b��wR��kd��E+����W>/�����Ʋ[��ՓH�˄�o��m������+2
�����(���ۙ5C4�hR�Kn�x��@�iqvF&V���9��~ ��}�<�����_����� �wu'��Շ�X`�(�友hh��[f�gk�9���@q&�9ʘ6���+EM��ɕ5��cAX}h,�[A>a�3�Vf�IŜM[$�1T��'L����1�D�ǂ���ew6�䨩���d�F���Dư�#�	��~äޛ_�:�E�(��˕?���vb�m�ø�U�	qx��Y��x?� Щ�&��w��LbNs�������c�z�;k��>1�n q�F��=O�K�,lK��(�+گ�[�z�sUt]���>���|��oD��	w�0cn~�&A3�\��\��fY��뒙)͈�dExQ�ii�9{�vINR�M�{^�\{��ڱ�\��#��$�z; <>v�Yk��8:�-��{`�0�	ȿ|̧BE�?9���7twĩ�K r_�#�A������~ǁ�#N#���FEV��/G?ݜZ;F���H�$���N��\��:�����
qSj�KP\�s�4jev\9��wW�y��Y�kSwmE/zi�'��ͅ�PR����~8���xÙ���3�<��-g���F�<��Y�g�b�du�`���
ထ�	#���elۆR��V�V��yr4�ث4�O��&�2������_���Y��Jxv��6Yz��9+R�v�TB��<�f|�yRq
�Mz)*:r�y���-�F_^�69�N�Lp!f���2��o�+EO�_\�IV�K.�$���l��O?#Ԉi9`�ca��IɿԵv5�c~Oi-н9�f���Y-9h��:�L9��0%)]��d�� �nj�3N3ї5�����Αpܭԥl��s];	�Q�
w��mm�%�Zs/�(��݋;i�[��+~��P���ң�&n��b��|��G5��E*��a�H{3ș��Ҵ��]��3�%!�l+���֔� 	)��W_����'T��Z�
�ӎӍ�9�������dX���IjTM��OSLʁ_����W�?�?蹐L�E��c�4A&�l���O�6�^��`g�81�{*װ�j�nl{�0L�'C乴傭��jճ�����)��E��1D2a|s{�)��g�[@��jM�`�Ȳ7�ٺߠȣ��?[��$���	�W&��Y��Υ����Z2n��y<D�hl�����@SW�QZ"��ݷJ�	~c��i��pBn)��֪Ą,Γ���^������O/;m���5���v)�5��o����9]̃e����&V(�����[~ŏ�/�S�D⻓+�W
G%z��B��W���*�L?4*�B��@͹U2�~I*��ER��^�Hޜ)�J�'D�Ҵ�D|�7�QRN�k%�<��/-�����7(Q*��Ф�6	�}�z-���X�!�r%q���� ��~�"��g&V��wH�92#
�.ŀ�/)����a*�EWf!2<�����`i�,�R85Y�.Y Z�M���<��(�fܽ�Jd���V]�-�S7���A��!�%���}	\*@�`Uڝr��z["0��`|F,4�U��&�79	�J�����Y�'�%� �5l���������}��EM��	�tŷX���$q~��nw�ugzќ3{@�ãm�m�5�71��\(������O�%�\k���#e'�\�n�y��a�J��jMhDUF ���MX2j��ߗe�!��f��QҬ�ڪa�"Ms�xz�_feO��v��h/c�'0�����4��t�@���=M�O��[���8!��Z{uks���C�5��&�߬�t��PK� Yi���|�K�r���b�H]�O��귗�s�����j�X���K��oS`N訮��,����R�iܡ�q��aI�Z[��,��-�A˄|��A�u TN�]���߹�X5�.��)�'wd\&]g�n�6�"��d�a	G 3���h/�����`�Oe�<�B�U2z͂0%�x�^F|�R��Zqxkb��.we+z�$!Pٖ�Ƈ� |l���nx��b�g�By�/C�Jz����]6�`�T�d-�c��J�6����z���G/�����`~��e�U|��NR�!W��������v��+6eBݺ.
E�h�&�.��o-�X��5�E�L�䐣��V�?���KgU��a��U���D�f���X���C  _	��9H=����J��eL��7��녋�d"[8m�ۊ�1tHr�Wj&��z}�KX8
p~1�73����٧�v~נUH�F&֙r��b�P6pz&%tA(ό*H���i^>��a�����.�E�j�ɾ?�*j�ZM��AS��?��҃�x���*��Az_�ӿ�Xh���'+`�m�B�܉�V$G7/�L���&?62�i���ZQ�J�\�y[7s��4	q�r�@�g^Ne��mK��n�Ք��>򕖶j��;L.VKD����>��ϡ�MǗ�R6���G�Q�Pe��& :J0�!���ua�2e�F��v�7yt������R;H7���{�V�uFPP@��,F�y��,�>
+
�Z̄Sb��� h�
�x����ҭ�ߞ�ut�ѿ*ԔIh���G��.��1�o�^�)��;��q�"�0w�&��Ǧ,�iUP�=��$Aؑ7Ķ-�U�_aĝ��N���f�&�XI^|Z#�U2.�>���D�ްe�&�������W�x���1u����L��X��2ҮdX��\��ik W�L�q��
D��̷��ó�B6E�кo��]��|7�B<�0� $�ճ��ٕZH�#�D{F��%�u]N��l|�i>{�I�޻z��h�֖⢧.�9;rGrJ|d���\�qz�W}��m7�\c9r��:��{ZI�ڐ;�α*3w���2ܙ�Y4&�-�TS,�Rg�����f�)�E��6�|�A�l�fOD�C��? =����'/��8�M�+����>>[�*�'�M�4��JԛD��� 	�Q+.Í��f�aߑ�b066}�(1�]�a����g}!����
b	k|�����ɷ��0m.���-�ϨJ��.Mo-�T����^W���L�ʺ&_�[$��ss]�(���2tE��xH����]����:0���׼&�!�y��������~(�L�6���4��h�`����WIʧd�8��9.w�-F	H�}�r�d@M���d�ѡ��2L�.�i�W����9=УBn�x�QԱ���I�%��1�P��� d�b4@����h�o2S0�:ҍ�${��'�T������-����o�
+�+"������xV��E�����榦i1.�Գ���?VD�i�]��͘� �1{x"���,@��7�7$'$=�o�����>{�%@����Z�jǋ�>�Νp5�H�Q򁛇��اFv�a����8�J�<�ͱ�P��L�F��ҷ�K��f��a�~	6���My��0�����OҪ4��:J�?#ebI���5�IM���� � ^R��u)��,sՏ"�gU]3�\��+����Q��״����	�و�\�8̇x�C;�E	�}L���G�!��$,�����|�M���6��S+�B�U�s�e����2�i�C�GT�h���"�M�p^���C���И4�{K�X�j9s�~6��JY�8��rS����J�AK���j�U�~��f ��
�nGZ"� f�*��?nq�+�E������VĶf�eDb�K��@Tb05\I�p $���f^��ٕ��s��2:6���"�%=���{�Q	,%U6�{�t�_�8$��/rԇ��!���˸7�ؐ��$0!�=գ�ї�V��v���H.]R��zl}s��t��k�54�C]G�~�ư�F�̯�*]' .��5�۬�[�ؠ^�C���_eSkX��Rq���a�5<SoC�V�K A���>�ۖj��h���ې�m�w7�6o��٦
�*��qվjڭ.X���.RΒ�Z���������*�p΋t��Y�r�����+/C�/��?$l.�R�6�1L�#�ګ m����k|����%jk���󳦜O9��*�\���{�ǯܡ��	�?-�;�#�=m<�*Ib��Xj��eZ���b���9
뎷]�J;�Y�����7iE��)�`��o
C�����/2�����6��^��Um��C�0����?3g`oZ�#_��f�?�����2h�=�
���>��?%�Rs�'d�Ь��}6i�Ә;�����{�4;>-���k�[��T
�E�U�M=d�/��0�h��[���#�.L|A������j~�o&<�_�%�^�n-���e�dݼ�DAW�p����9�iP�TB�w��x3�Ȼ����O��\D�=�j�ԅ�'��sȥ����?�/��hIW�8���z�k�G��ʞ� t����oH��Ŋ�'+n�z�����v���f��/�d=�nE#��?WH��m�EI��7��V&�;(.������08���X9;�k�?�a:S��/���7vQ���_�'���S�a?��g��W+],�gHD��/}$�xJ�2.�YYL�� �7�E�p�ܵ7:%��FUr>lR
P����9y��ZB�wF9N�����S�u�7��# ��Io��/o������(�ε;rx�D�
)�2����l>�c-{����Xm�	����ʕ�;�\�b�r�ԭ���-셎��_�D���l�B�J�E�I���S�g�ö#���#^N����y�t��8�W����~aNE�44��zUj�vo��g�x��zhFl��\k��s�G�B�驴]Ο��o���@uO��r����Y�,�G��f;�a���N���C�IՎ�����y�\�{8����joΰA荭=x
���%-���a�*�����L~	�Y����a���`q\M�?�	:q$~Y;՚�_\�j���_�x�M��;s㥥O?sƦE�׊�G��6���(�vW��.f~@G8�N�����Ml�	{�N>y�c�6V3��	]"�J�M�D*���ʌ�6`Yv]X3�r�`OcZ*�������?�@w�d�M^7<s�$�u�f~m�N�'���$�����$���0f&.0��$&��(b�FV�&��[Գ{ԍ��ʒ�N��9x�X� �+�7ޏ�*\��6��6�Ԝ~6�C���q͉N���X#c�kt-0gK��H������*M����N��8����:�k���{�z=�H�_����(xD�v,vDY'�٤Y�0�q���ìMY�֕z�d�12�m�'9��9qy��+�[�m�����w�#�����j�妁0mg�
�BBh��U�~�������L'L����A�X-,��$�F����Jy�%�$I�`cv��/6��)?;4�{li�[�c+�q+�.�9�q?Ӯ��m��8����r�@����YH���O�^���
�S���W{o��! PiD�)Z�Tŀ��:t���,�/i���O�Tٲ��(��x��� "|�_�}����j��mG��)�j!A3�=�Tr�Q��כ���:��SޙRp5����4\I��ǅ8��k�k�(kS��Zw��`v��|������? �M�i����H�@�V�O/���i�X-�Mֱ3�R�$�	�|��G�m>dj��<�N�q]���zZ-�roI�Zo�ưWꬃ�Z7
��gwhlD���v��� ����y<�aU��J/�YC���vݓrH݋֢$���?~�4Sʚ�f��	�����F�A�9�|���i��C95qS��q$��qR�&�\�E��ei�o���Or0�ǐ�[�E�?�/�rQ�ÿ~�v���ٶ�M»q�v��i��W��V�x��o��Y�q���q���O<�%&���p�[j���[�*"룰9�*�s��0��i��7�'�h�r�m����n�B�ҡ��c�l���?*��F��*�9TX6��I[�bc!�F'�H������B �B<���R�]Gr�$3�~=�p"2á���[>ɠYi��r?�_����m��%�Հ^͹�����#���A�x{�'�OJ<M��b،L�����jxo�\Q͆E�Lg㣜3���4��ܻǍbC/\x'�k.*	�`�4} �!�����̳�A7��TB�y�7���S$o �ڌ��P}����Ӛ�;��e�v0�C��FV��NŢ�0��qCHn=�u	��b`]�qa��k;'ݽ�ʹ+�~������s���W'p^룬\��@,��+ͰW5�o�x���W��*��� $B�p���+U���	��zxnP�!�Q��a֗{ِ���!�Ǐ��(Ӹ��Ab3W�a���ju�!*�̩F�P����3^>���;"�l[�|���t�Bl�	����������]Ш6l�i��'�O�d�x�{��-��dP�l�����q�{{�̓$g����A	�%��B�v��;vw�������o�2b��5,m4i�Il��N�V*UT�؉-�R����Δ9����0�����8�f��sޛ�2�x4���dQ�&JNXɠQ��|8OQ��x�Ǖ��u�UM5Ȫ��k�̛P��;P��AꜴ�}�E���Icx��s'bo�#v�1~R>��l#M��fx�|ظ�\ �I*C�hi��7'�60�>���֕Q��02+&�)�~
�`�xF�;B1�fj��'�=�V����%�e�h�GP���šBC�C�n�F1��QZw%�[�'1�e���@��i��%q����3��V�5M�~`�،�=8��-�K��������n�r2'I��kW���3�O&}��NU��+zW[�篦������"`&y��G>�*��]a��iY��'�;^���H�v�$��;
t1;�˲���3�U��R8�?���J��E�]���ME�kh�㶨ǅ�2��ģ���G7�_���_ڃ����=��OM�]gm`c��q-��@̗�˿M�q.$�k��~̳f��Z�t(ʛf��5��x���SU����nթ�tU�v3$��}0;M�V �������:��?p���+'�⮿��(����A�,Z�½����}�̲�"��4� R�ȹ:mo��kG�Pg<5����Y�{�� (h�KЍ@�6ĭ_ �ט1�P��T���&007���gv�J�����.3�P�>�IX����G_�k�U�,���ِ!�y0=�N~�Vjn7#g�M��96���R�������<��t��3���U� �gF�V� e�W9I"�tF *�*�zR��LuL~��>�j���néƔ���^'�!�נ�{��ofxb��_~��7z�8śm���R�a=IO�~17���NR*�\���a��w�*�7�R�v��Ăo��1�PiN�P\���Yn@G���bw���r��;T]��f��Q�.�ϝ������y��l6��=x�����|�ϫs�{T�fS-U��dR#��Z	_K�5�B2��5�^���R^�s̃mjM����$�d��]��;L�;]Tn�<B��|"G@�M�Y���T�1�R��[�}ÿ�/B�Ħ��g�{i� Y�m�"�:���WE� d���"O��r ^؞�C��Z�zk��H��nU|���<�h6<��*|�gJ��V�~*�?B!ُ�_�A�:�A��>�1��k�||Q���ˌ���D��V�e2��,يc[�R���{��~L���`�ۃ͂f��4�6�3[n�j��(��@��'0dF�%qc�e1F�BNfĞ(����ϰ��.�&����7���3ѿ���<i��N�ɘ�wjN7zwi.��V�����R�/�&����_J���t�>j����L�~�9�����_}��i�%΅\���	:]�?ؘ�Ծ��M6S�S�YTT|��IӨ�`�$o~t��ڶ�W��3����`+�u� !{�'�Hq���<�������l��������C�GF���.�\%��0��5ў�R<�V�]o9X���5�z9%!?��+sN��+n�������-ǒ���7�o���]�>���\�����n�#�|��%����p ��H����]�ĵ�]6�$��I����텙��n໏������@<�|��	�I��+�
����V�Y��#�O�뇺	�*��c�s�J�d؛�l�$�"D�X�d�s_>s ��@zq��_Bp� �JWS���Z#�HPµ��	w$�m H_i	����N��5 Z6:���EQ�!��hN�~�x4�;��p"�2�=4C��vҲ?����T���Q ৴�k!Z�d4$��}�7(�����X�؂ #)�V
�.ތ/Դ1�
}�bq��WAeB�ʅ˽_��_�7
�����/깹��5���iHm�V)"�0�ai�X�]@�/�:�����2SC���Ry�I��?*� V ��(�[�e�2�\���n�O�Ώ|���( z��1n�Q�:-?�,�:�z?)�w��.M0���+ڒ�a�T} s�Y��.��t���"�Ba<�C{��D��%P!Gi\�sm�����"� V�Q쩋D�7L�d�kU��2��
��?����(j��F6 �]5W�\�X�W��Kn�:2N����U�2.L�_��j�w�ʊ�J*e#t�w��$�KS�sL��e�u׳G��CV�cC5o�9=��1ç�+�r��2�Z"��wo���g�ՀK�i}K�A�T���ր��Ũw���_327���Z>��+�޴�p�x7��%~Dc�2OO��;C������D��՘#�{�Y���W�@/��Io�40x]�T�����n4<J�֓�4?/_T��:wP*c���2��OPj<$�q�Z�����O���Qp~�,��33��%Oɮ�Q�0}E�m��$D�.�\���C$޵O(v��	�F�]�BJOOZ�R���춉\�*:��B��1x޴���~�ݵ�N�,4q�қ�'�!��_
�Hy�H3�%�~�D�������+9�	�UR���7@���� r��ˬ2�\���oJ��9�ظJ�����۰h�GS��פql.�Vg�3���[C����i�9�-	�Ήj�u-Wvm+
���� c��Уw5��?g��M��8X���(Ĝ�!΁rd]�� z�]�iN['�w���1�r1s���-H�'˻�l��v��1𳣔�g&(�A�
��WYB�@��|�pj��ғ��*�%W�%ʑȎ�1Ĺc�s���o���:_�IS�T_����?�7�	�l$�*��E����o���	-�^�!jj��/C�=ڐ�Uk
�ݚ�7�·��`J��n���nCF�`J�;8K�܈��8��v���
W9���SX��3~�+hu2�W�@s�ö�KGs��9��OjV���R@�#�=3���0#��c�Rn���O�4�^M�坮��î�U�.���hS��ٝ@�g��IM�_^����Q���;�z�7N�����E����[��ؼ7sS�:U̬�$�]�Dq�S:nf˽�+�~�����g�ox��F�!;��͚&�}}Yj4����S2~1L!&)��qVqaϪ�.�Y���ka�V�x�\�k��)@��J٤�/b�;�-����U��>�`���
'�4H���
a��ܯ$;3���|�]y��'���	Z~x�t��k���.]�����{^���%�+�G	w�R�xM�fPEP;q�*íԍ	�Nn(!`U�L�,���ާ=�0j�Z��2<i��>U���R�k��Fv���e��2�Hx���?i���D#�6����	$�%�]^�/P�����*c��C���KzL\���^v�}����G�/��,�_4V�`�ٚ��AURې:/��>���B]~�J��Cg���¬J�TN�/��4Ĕ����X7x� ���\��i3������<�����8�
�C�s_���d��u�d\$��ʯY�n�
w���n"�߇��HX�%�#84Ճ>.:O���`���L��&�+�S��2"W|LM�@�ٿ�^dteV�D�����Ї�G�,�&�BT��W9�����j�����쮩���5�f��Xd(�4�KNp�S�$���~X��`ʗ����>��H0C��m�}!�,��A�L���c��b}䓘�R`W� �q����`�BF�����F���*���e�ֳ.�7��`H���~!D J8.Mъ����3N5�a����(E���gO^�����T=����m��W�	�=$Ƶ�R�����n������,�9��� l3��H ��\�*�E�E�W%�^Mzz��(+G�������r�}��l���#���o��mH�n�zA��I^3?��� }��T�Yh�0�f꼦Y��X�������������^�
%�}_�?
I�L���"���_BQ�����<�u��8�haĝ�Q�����ۀ����ZD�HF��%1�M�wwrx/H�v����*󓤶;>��^�,�����E�������@�Ng�P�_m���l�"����-��׮�r}��ˋ�*�������B^����L���6�;�ULsăxV3�x��$���7�,L_��Scm�ᯩ���e�W���#�hg{�HBW?�+�)�A�[���A� �`����	��` q}t|��	3���B��P�>��wo_���V{_����ORij!ḵw@�uC�	mǛ��d�˓�1,��`�~X_���y	1\�d�� 8�9o�hs~�������iD &CoS|(����S�vm��]���[��st2�����2��lE	��~&D�F���{�@i�Xf���Gt<��y%�-|�}�4%a���a���:;B}�sFpl���$v�p���7t�u���=_�@������F=�Y��ST����-�����=�Ƥ�q��I�F�rd�$�@.�k�0@H�}FC�7��t��B)h����9gq$?��Y'\`�f�PgoC���l��uN5�P�6���-b�@��m����W��X���<TFa��Bk|��}7�c��g�zzy�[Dp ���f~�������nY1&8	ܛ\��5�ǆcz>Ft'���W��'�ļg.xM������<�b�x���uJH3���V���� �ԯ��ϴB�U���;z���ϊ��`���ϋ�<@DE�Wh(�!�����H�6���r��������5�,����~�����"��^�� �5bӐ�:�Ûl����u	�Ӫ�@�I�lۡ�%��y/(��9w���P�5_A�P�[�,��i�
<x��k�'�&�%+F(Kِ�����J(�wL�<�hҤ:<�P��W��<J[�@X�������k��P#Bd1O���M��ް���dx��}���9& ��RH��`��+%6�r����zh4V������U鑯F2lq �P%����LR����.��e�C�ZfV;MB������.yM�ɽ�J��e���TJK䂪V)���*��'�hJ�S��8�i��&�ϕ�����![�F	�{�p�E!������f�Øz�C�����k���ε.P��~Q� ��]�e�#���Rg�%4�%�;���^��Kܩ�(i��M����Y0����t����j�;��E/�K{��齖�X�H'OGE�	}��p0��!a�i�c"�Nm*���A�t�ߟ(j�js&'V��5�d��(�/#���dc�W��ɲ�8F;��uCʷ��{�pn�v�����*�/��M��yK3����+Q�`k�=��:pK'�#� ��q�����#�D�u�]a�P���J03�2�;G#V"�؄���w��+���I7���P�����H����G�;�OP"'�H�1(K��0O�\����
�oH�I_�n,��\�Z;�Hȫgg�a�]٧埤lXN����}1�����y@�ؤY�H=$�o@�<�]�A���Ps�P6Q� Qf?�6���ꂪ(BBX�FS+�_�^8�*%`F���}+���'��m
($�2�g���IpT=�K9�;�7R�̵Y�$\����k`*� 8T�S `����-���WcA
1���՜�����o���u�����S'�N`��љb��sȊ�_�h�#�:��E��_�Z���q����Җw ����z1�UjN?sq��W���7\I񤬅%�9m��q�x$��o��-똌�C6���c?EP}F�$I>	�(/?����E4�]�p�2�	��iq���������4�����WN��dk���g,�&��+ICx�cB��7�+�h �P��r�%��m0�������d���7z-k����3^r���xz��kO�6�{�@�bF�oÊ�g�osR�W���f�2
�%��=�X��v��d�&����Ψ9�|M�6��թ�N���Q����?��w^r��:�WQ�+î����U�(�p���!��r�ێ�5
*rqb�=t�a��\��"j�?H�A��8�K̳m��y/��m��B�pv]���9����rhx2�m��
������ȉߓ�׮�`�ƙ����}˫�����D��zj�w��!j���?꟭�/����N*a*�M��o��rGIK�El��`�/>4�0,���Z!�?��b!�������d�Ω�W&
CM�Q�ߕAJ���g��)���[�|TV��s�x��>g���<�>Op��j��� K�&̌ w��ͽ7�	�]�� n�Yȹ���D��,���
�׉X����iW����G�ߤFt�+A��I����v����(���:���L��8�����/�":t���ʗ��NBZN�@^�����r�5��i�Gk\�8�K4&�?�U�.�	�кi^���C��t�R�&�͙s2��$�fZ(2#�����r���;���tWKH[2��H>���[����d���g��b"�����ԸZU�B��x�%2���]�mL�
&[��� �y"�C�6�-�c�&@b}*�6�$��T�+F n47ظ���G��k
\y�G��aJ6�nz�wWÔUk��l��/���:��f?8go9���$$�9n�������N��B�ތ��3p����/������5�,;�x�VfӮ3��!U`nT�"�"	a�N���@W�ݓ�=�b�x\C�E���{��P���>s��瘫!���6��!ޣڌ�8P��=ͼo�5�>�"}����i�mYB���Eq&#-����X}�9��G�_CT��"�=��Ix���5ǡ'׵�,!��m*���E���bC���/=��'�l���K���`9L�M�+���r9�I�@��?@�a�z��n���[�Ku��WS"2B!
�X
V�dq�O� �D����MJ~0����&�� 2���-:,'�՘�a�U�j<J���/��{�T �{~�<�Y���8{��mM��K���8�Wpn0��D0bف/J+67�br��dn���L��W�����rϠ�7^t� �28k�E2O X�<���R��dg̔vd�Q��϶�R������	f¯,SYU�L���^jg��~Wa���'I��Cֆ�MX�Fl��amD�E'�L���D�7��ݲ%����U%d�*G]�\�	�q����!���j��	Y��s&U�)�h!�o22�~�u3��|,�i�W�-8�����㥬�3ҵ ����!v;�X?C"����hsn�O� +�Л�^G[��eԦު0�j��b�t�Ču���0Gy�\q������{�J��Sr7 w�Wk���W�mS��TʡՁ�w���aUtz�p9O��[:';/կS��\�qmk'B��U�8�#]2�t6��H*�$���fe�m�Ê��Ӂ�����]���/�y�P�j��GD��2���n���HH���O	�!H���.��#���M��>`7ӈ-�hwL���玊�*��P|(R���.z��������#�1��
��pTq�Q�Eoh��@��$O����=�P��x�j�|������8r-���]4҈J�9�:�37ؕ�e��)/?i-S	��g�xJ(�m�"��b�QL��z%��y�ח�ƚT�3��l ��mi�����*��4	zd�\+��T���S\3��$b1|=��d�ަ;���������7���wfk�=;��ͅ4�E�]�� �wD5�H] �mͳ�<�]��bb���JX��v�B�{_��n	[�R��ۡi���I�&p	g)<K����}�b�%�؊�@w��VMl��wyg)�G��mz+�
�JD)_b���������z�JL���o[h�p� W�U��c�R�y~D�egM=����`���I���wc2)��~˜[k���#�8Q\ᑹ������
�>8%���H=r*�s�O%dwxcy�*5p&�>����;�؃�Y��E�^D�5�k��yt;�9/�y���&��6\�8.Lr��\v\�n�͓��O��N���& �����b!9��+��<,���_���~�P�)]%��;�%.4ff���Z�~���&�ܗ�:j�^�'�K�g������/J��OYX�Ϻ[5���_�#E�p`ʾ��4�Ųl⾕~����O�:<���L�`7��y7�>���4���l����6�@���e��m����*���bV�)	s���2�E�nA2O�Jn}u�$3��{y��X\���8[��[t�/�y��5����  [��5=��
Z~+�Dٕ�H��ʑ�W�`��{�� �-cU�X�I�["��6e���J6c��'�����X�t�NfUe��s��_��_�O��%���J\�	�����/#�D��\�]�tzx>~��� )#<Ac�\̼CW!\��f���u�E�Y>ײ�~v��&�u_�&꩝7�K��'���_�l��IF����辻�0�A�୽��J�:g%��}I��o�5���J���:��#�]��Κ,R�%��>I���W�Tr �B@�!t���j���ՉIٞgڼ�5���4 HM������ow�����\����[L�Dߡ�%��#�sS��(��a�8�t0�l�r-��l/����Mu��&����Kp'%Y`s�t�t�I����X��Hs\h)z�|�ݰ���[Jxa2�rI�q��f�E0���ѵ�+vd]r���vI���	��HqE�)S���#��!S$�}��yj�r�4T�/pË%������)l�^Cřu27<�8��}d,���w*M�^���t��z:>����·$	b�7��_�ڐ4���`���6��M���ZZ��*�._:��O-Hj�,���P��޿�\�`���
�������+�Y�"�ݢ���*�z�Er���e�Wr�÷�����B��
��8���rO��;7�2af���ˢ�i�/�ͅ���\5�л�1����YJE��~2�ج�0�
Vm�:L� �tmˤXRa�?ڋ�n�y�#79`QC������#�c���P��9>C���ଁ��n��Q�;,�rWI�Ҷ&��;~�Dϼ��P���w�̀?�+]�Gܺv�_���&i�6�,�7f�u�[~��|�y>�Y�d�n9��#�0�,u���0H�Ab`�K�X�I�	�w&~m�~7��%)�m�3+�Q����	��o�̘y�K�nL�uj��qR�,Sg�z���M�n�_�:�\YX�͜��J�H����M3��[ӎ������j=v NFX��!�}n�]x׏F�`ס&��к+2��0l��H�,��!���X�}ns�F�U�p�`�/�x~ �� :r/M��*2E���2�)� ����-��9��$�[�z>�����̮���EA~�L�FCAo��m��nGA� 1�+�\������}7 c`P����jU�։Y/�.�(��}��òx�w d���q��Nnvw_��_ȱ��]�	���jX���a��Ϯy��i�i;�)TӁ]����s1�6��\��L�?��8b%m�p≇�*B�B�ɔ��˃���9���sGAբ*�ZG��7�f�����X�6�Ʃ��z^	=�������&�I
����^S��n�9J�Rx(�����YX�S`A�uԿ"�u�`V���������u��V�x��7�����?�~lc�����o#2Bk�k�>��Rg��{����㚨;�pe�=�+x��u՚�����
?�S�"�P�����%�	~NO���uɓφz]r�s�%��;����ؿ� ��'�*z\C0̞��ױ�%�5��`?bh1� usl�c��v�x���Nq�n�G�������[��S#�\����מ�w�5QDU�b�k�B�����[��K���%�6x�\��i>�}�@Q4���3(�� ̟�|�U�x��6z<�ő��W+�Hgh��!�]���mIZ�ݎ��ڠ��yuؚ�#nt8c��}\<PZr9{^��^�ؚ���#�۽67��n��q���������h�9� Z��y�Z��r����$`i˒�jfWX��'|\�%��5�bM�ĺ�Y���������Є� ����(@�����r!�1[5���!GÊ� #ފP�E�Hʕ���g������g|��5�3F�BA�$gۗ�=?V���L/�"�2D�U�^�rh�ō�X�O����q~�e���8'���ϱ�^�L��ǧ0P��D���OD���rB���\����I�J�ҟCxf��o��C��>�Pu|��irw-0-+�������H�G�l���V�(- �GgX��y揶Ed$ ��s��}mr���N�RMZ(���n���_�^-�� �=*Q���3R爽/�U�\TXa��A�)��ڽ�}�3�^X�lb�r 6+
R��M�,�ՅD��%W�S��2�r,�<��0����8�ޫ��Hʚ��E��0�ֆ"�Nx���Ft/Rvv�%a~
�"�$D�L�f�����y.>�;8pq��Gw�=b�{`Jߕ�e��;�~��,��� �	�����+7I��D�>�(�MU�Z; ����~��nR�f��Vݺɭ�bˎUwʆr�3��ʭ����
v��ཹސ�B�b��:R|v�<�]5��g���m�/ k�P��b��||q3KY�=��|y��GOrZ��]���sU�a�����r���9��w�8��(�6�a]ͤw�C1�#p'�dw�0�S�¥$sǣ����j÷x��PX$9̧�E��L6X��Ti���ӊ�������.1$n���́ �\�����08��uU��}��ȕ�M�=�GC=�Hɠ�����w��N����ߙ3����<ƯN))�r�����qzIXI��	�����S�]j��3�^g��#�[!U����}��m��B��i����]j�MJkf��Ӹؗ%#��O�X��k���!���iYX�>��<�K�,1�k�gD�:�S$�`��mOڇ���h���!�qc�ÇBrȚ���t��w�cy��j�q�ڱ��2���N�q/�׸�2C�U��׾mµ*����9��p�"��V�L�����0b3v�����.Ռ&��wa]�Ȣh��ޕYuxԭ��L���L�W����c��6�g u\O��'k�7D�dRF������Z�/d	��z��BN�Ǝ�H��g� 2���m���Z�h�%���
[/p�s�A��b/K�Q��)�U�J ���Ψ�b�Ӄr��+��������Z���i`�D`������c0�~=�㭊��o+��?��mĐ��e�`͐�66��ևw�Tz�&i�@�F����V�#�^el�R����GF�,�+>��d`�H�)�5��^Ɂձ�S�*�푫\qM�t�8?��D���R�[��ٻZ���Gl�>�{k�L�%��I��ଃ�Co�
Q4�=n_�X�_7�h�� t�!4�f��e��0t�|�Z��Wa�����G���^]���g�)-��"��0��{���g�eٳ=v��H1H��`�♎M�Af������kFz��X�ٮ.�ݕv�\�]��&�Cm~�;bh���T+f���>^FY�8)ԶX^n�v�osǩ�]@��
��MkU0kG�/�l��K�w�)���y�g�8�ܯxG�|C�3���+� ڨK�)�n[���Ch1��JMTAL�<�bbFSP�p�W ��Zn��^pQu;��/r��T�zdTp��^E]x=G[���տ�+��;���\+��lB
�������ô��ŋ�(m��/ݬ��n�r����ݝ� �/V5����B$V�7	7TMe&�J�lr�났g���s�9�+�T[���4�[�h��U6���hI�nc�<'�m���J��#�%yn�cC�<��6*�nz�5�>\��c�AF>����n5 ��Kv�6����>3�љ}z�LG��e_�U|�&De>�����֊$��X��������E�s�Ҁ���8aQI��>�U�O�_4Ok�s�m��'��3s���3Bܚ���ık�x�^t�؈XO(N��DSa���D\�!�L"
u��Ǭ�;���Ct2��R^A�kj�7�8�������j�:*�����o]���~�m��`#�;��6��`>��3ê�})�0����x��#3�{~�?�G"څ{H�j`�ҭb��y�V���;4"нQ�Wn�Z��@��k�9Bi���y`�l�yR]9��L�)3�u<�ݪq4�M#����
@����mcx�����������?����P�d.�����T/�٣[y�ƭA�-(��Z1��=��!�R�H�����3ȩ�E�.�4 -���ֱ�7��VXaQ\y0 �|��
�ye�f�x����"�{��yܒ����c��A�D >��	0Cك���pRܛwnF>O�I���s�.�s�~c�k\b #��|����d���, oi
ʪ\�L�������%=��a�ה��rQ��m�D�E��Z��fl��h�STM���Ec������k�b���9�P�RFW2Q��7���o��|���*�r�/Elt�ZL>����ڢq���r�`���ϸ�����Y��%Wu�1�D;����Z�F���� ��x�os�U�ϯ}¡�@��=^fM�'$`�׻+��VG6��pqe/B��r�`af�^C��H.٣�b����թH�Tj��,���V��~b<%i�^�;F1�a��(��ld�Eh���'d1X7e%"����S���\wAY1�	���Ez��z�Ԇ!'GYR�{9u55i���.ְ&�Xm��(n���ZG"vb?��y�z�����\Ρ���z}��8��:8<�Ўd�X��Ţ6��
�Z��z&^Lא�g*㦷'jIt	�<d�i$׃�##��v鶿�N�k�gNj�Z3�7����ID\�< *��J%�{�OB"P�<�̍Kr���@q彛�,���m8�=���P�U�e� 5Q[�ގp)�����߿�\�'������0�|�+`۷��X�8�� uX��z�/TV&�����<���ԫ�#�d�K��ݵp���������XJ���M�.ǖu%�EM��ӥ��M�v� K &�Gh1�p�7�5��)z�2ze10D��!`��W�������Tfq�)�Z�`ٿ)�:8>��!�k7��M �� �%-p������ӑtk#L�~!b2�W����FQ����\�*�zg����H:��tw���A��H�JX�:�×�a��D쾽I!g.�����1ʑ�<����s��m��S;
��-�:�=�B6�8c��������^E
�\��B�p%��[�pѦxb� ���HC��&0�R{/<%�J�����(��Az��Z�f��u���&ؿ?F���o�w�D4�a��_�d+[B��Q�|�6���(k7L10�w�ܣ�-�+̵m�F����]�̀���ܨ�3�j�e�o�@�\_�h-�%���Ĉx�{�_��mUي�kD@l�5��F�#ۓ�0D��[��2�(T�z04�n��h�HkK�j^����>���A@��o��h�g����@:�8���^Ŗ)�r���'6�ɗz,����)K��c�F�� H���,��|jFg��@B5]��T.�0�sv}��i�m��q���-�ǜi�C5�?����+<L����,�����W�`h�������Q3��O*5�����iBK������\蠶�$�:b<��t1&l|$;��=$�>�,���@��YM�\,t;�Y:bȢ�È�۽��i�xX
*R�҃�£`Sh1��d)=?-PM�9�&V� ���@��̣9P��P������^eͳL���#圴�HY�Y
��#&�T��8i<� �Ṫ콷'�@z�u�#i��{U�`��Yh ���c�y��]��~�.�N���a���Vܫ~Z��~]*�톡��X�W� Ar��%��I+
!
���P�������tQ�4&_h�ܜ��W1]�.���4�����9!f���x�ӈ����?hJ�(��G�+bp	0&���$��	�~EFhX���� ��v�~$��Mk��ts������L���^d�m˩��AL�Xnąp�Ō��d���Mџ0�2&�
�)25��!?�1j��;2A^wﱛ��F�'&I>8������O����,�t�4�e����c���\�n�Yd@'#�� }�)�P�ҹOUb�#�긶���5�<���&7��qP-�}����K�ĩ���pՇ�%�̤pR���W��e\RW �&w�PW��J�X��L��}���:\�qV��I�,8��yX�Q�!����ad9�����$���u'z�MX���7]7wk,����.��/��~u>1�O�4�w�V`��]
r��ڡ��Hbt����l�X�%������7�>˙$�v�A�v#0���rL���h{F�!y_�W|����3�����p�0�K�s|`���������������}e���hR����*2k��u!�aTr
���O�bn+W=t�Q���3���x�ץɪM�9?� R^�s�LfX{8(:t���8;wHdw��'gW��]q^�����&�wW�:<8��T�@[�	E%�l�:/1�"��.��6�UI�!N�m�YR9/�:���9O�/���A�#��t(��3��t'&��Yх�wu�k��<<<Q̈́�A%; �	o�gE��"�c��į@�&�1Ͽ{m*EX�ϱ/�}56&��RE] �>,��X�lYE�V�JU5�nm�q�W�%=�XPT�!G�)C���[��@2�Eȼ(շ?��mg��V;�: v>Ofq?�SLX|D���7��;i���uR��`Z�X�#���!+�s�pIkf�{UJו0�꼽�F�ݶ��J�P,	�#��$�&ج]q��O��s!�����ir�K�j�fr8�z'�>9����1�a��4��� �V.s�҂}����0p�$�~А���(�R��|��8_)���T����M���r� xy��*Ɯ�8a�'�g��@v#�k��|�֓��^��US�N����yϲ����dw �n�����+�E�����5�:oᵞ�N`S���-�F܀�JH��$������aF[??(���ZX�ۋB�cЦڼ*
���<a�m���r��y�,;n�#��9b�����*[�p���I�&��:bHӰ�q5C������^9i�i��Vw��j)�YK�6������6.��z�˯0���h2����P)Rk'�Y6����X��$�.2/ה��fO�x� W�	3
Ė���<F�xD{Ckَlw\�琟҂©@!�/�Z��*'aL�

Ş(��{\�>m�:�)*6j#)�^�sT����U�^_�MBxzƼit�8�y~R��ı���<���A12B�vrb@� �O�W���>�2V�����^�B7E��,��B8�/�T�#��)���]�o֐��H�v�1��	a~B��0\:*��FU�<���:�����;#���{_rM ���B�����ϯ�!	��j	���-\�x�A&����M򝲯_����%6�3�e�=��EC�!�����S�o���ԡĘ
a�J�<a�ɉ]`]�Z�!�huՍN�WJ�$ϳ\��?�F��&:9� �ձ��^ye���sdL�	N����L��x?~kkig�n&r7�/|����������L�
�3T�ZS��'�D�V�=3_|]�h�׋,[I1 �c�J3	���D�'��b�m7�K��?!�b+��E��ѷx˻��72�!�J��>��E�.9^=�j���uր{U:�K�/Kt��1Ӊ����s�n]2��SOb����'6Z��쌙�0��k����1���9|���6	M��
�#ZGvw�l�x�ܬ����߹��#��I��zX[*:!� �����4���Q��eܤ�C7�[&P��7�Ԧ�D��y:���N��6��䣓ȗ�Z;����.�Q����"��Om��P�0�h��2�!�:mg׍	fц5f����G��?�zo"Ǿܟ�H���6ɻQG�Z�ԓa$�wDxZ��i!7Q�#C�>|I����'��D�����DP{Wҍ� ��(B�e*~Q�`=>�ۀ*���$;�g�4^Gg���.0�<p�d���t�Lx�G�j�Ll��"�Gk0I%�!FJrl}��,O�'��]A�����<�	xbQe��#*O�n�!���?�ԓ�� 0(:�DY@�1��)Q�'֩��*�*�x��Sp��<�դL����βM8Ihi	��˧E6x�%"��O�C��Y�_��4����5����E��NY�c�Rv"v�&�����+��W{��~��Z��s�X��Β�x"�m���36����j�L ok<�h����:�8�]nn�f�᪁N�l)T�|�2!uś ��}Hsv���� ep)���<��J���T��|�-:��6�$<V/$"�����x&,t����cg�B\��_y�x�e�P�ۺ�կX����e���5�g]"��u6�j9���/����y��O�Q4�AM�p<�j:<�t�o��t~�~����.Y-�'��oN�K_�ǑKf�V2wl�Q5�e����Ơ*醿ө_a58�]���nSL,ݧ
B/�&U�qE".p�Y$�=Ԥ���+��p��u���{䢐\�Oз�M=�Z%8�4�ʽ=��f �"5��5{�eg
�Y1�ݓ���֛T�NX(�%(��{���Lq!-$;f��(���Ho|��G9��j|��m��4䛴4J:h1���C�åχ)'�Ӎ̼l��i�Fa����71�L��x&��Ǡ�������+6z��Z������a���X�琋X48S�u)	��ιH���gl���j�+��Sm@���=�稦���Ф�#!��c�Πݯ�"l@/c�&&�W�����,vx}��զ1�Bp �X�G���8$�$��(&�@瓿U#hWI?p��MX���ε��~����t��*���9���2uo��*�e?�d{�/|9;pz�cK,j�c�\�=�j��Ь����!<�몿�m'�K�P˩��d�耳/}Wᅖ�d�|�r���XѬ6��Y��wk��u�B^D���,E��%x�/u�>;��6֋�y4��t{r/VA�n���֯��V�o���g{m�C�����˰g�D�,y���$׉�Ft�М9يh���=N/1�ɝ����l��&o�m���h�V<��g�-��#�ֆ~,h���4��9���Ÿ�����_���&|�2�p�[]���,�& ax�G��e0��xf6^���%6.(��i8��S_5�O����@Ş�cXv��1D�6�k�&��9��	�_
��?UD�,@�4�!'��v��'Ƴ�¯����Ss{s���Nl�M�b?)��F\�oČ�����0�$;��۸��u�`����J=� =���{��C�w� ��`e0�?�	��@}8��.���I�)P��A�A�$z��h����������<�{�W�Izo����RsuP��^��$�W��A4P|�����}�pfzP�Y4)�Vq����{�Z!�ݠ&>���N���G����$S?�t�/J����'��_ �F�.��(��9��m��0��sP`�[��Y�Y����3D�G�!��%ܞ�7�a���H�R�~���xl�k�8�]�Ð�.����WFze�U��?;�gY�ޔ�q�3D�).3[���tw�oj�#��kk	�ݿA��*�ŏ�G"Ma��aD�A9��ƥ����l7���=*5��+�) �dy�h+�-2�fw�a7��Mt��t9���	'���MI�y����zWx5���ρ ;��+7!�%�p#,pҮ�
G�:D~�J�]�VM>&��zyy�����f�چC�P�_غ��4�b-Էʗ*�]�=
%�����b�ς�_�N#��{�����$�G�s�<�Q�x�^���p�����x|h���wm�2���q���c�8�����a;$F�F[r�V|@I�Q{�Pm�z�׀#������[�I}�*�gW���w��;����$.��dJ'jԙ#�<�m3����O�x��+s����y�YR��G�ѿ�l࢏��jw��i�X��n0��i�V-����Ҷ���|��m�GN7$�ZWZ4�s�z;���f��rM$M'�&���?�$�~n~��G�loO�ad�$��l���~����>����y�0��B�����	TO]�OAd���>d�$��ߛ�,�@��ek �y�r�o�I䰘C��I�7 ���\+6N��KU�B%������?g,�j2������AR,��L�i�H�i�&_�r���J�%,�BÌ�s%��^~5�	
ܠV�Qm�<�Q�F�s{Bh+��.���1�Y>�y�>��A����z���,o
W�����x�����T�ܱ�Ep�.%�s��F��s}|:�Q�-:RM~%��֕��n��}�Յ��9+_�v���L�Ȣ��$&�a��`��ey�d +�M�uZO������\�*�#��7j�&pٸ��=��e��J�s�{0�� �t;�D�&�xXp�o)��l�B�(�4�P�3����3Q�u_[��h�X�4�%}Մ���qf5��ǣ�.3��?A�|�p�(�OQ��(��m�Z׎J�V����L~�΁?G��pk ̥QI�F��{:,!1�(���A�h�2�h�vdW�����8���'��}Z,�ܯ>�@C���n�ÄS!�>}��v�K)|m�Wu�ηg�y%��HcL]�W�C!W3o-��y(��#��>�[z.��lpP�C�d�o�f��wy������WcK�eZ���	�GL��Wa�
��2Č��0��/m��L�عOq�j d�4�u�ȺJZĻ$i�G���ig��ډA�Ö�i�q�Eb~�z���kܕ�&�@�%/���|����>��0,�X�ۘ>��m����1Z.I�:�ٝ�%'�&tH,5ߘ�=�3 pP���
����4���jt��mO��v�� OXk�%�j1e*�p����b[���<~�c�';��2��:�U��L�6@'ՙ�)���D/U�Ր����|:����*�r�����%�]��̞��ۅC�_�q��������־ �Tc8�O|>�a��1|h�6 4�a����
���"���O�g��CSk�z\S�:����d*�~oМ���iFZ�l�{��NE\�+˥ �#4����c��c<�1��#�W�Q*1������nY;�(2gH� �C��(ː׸�O�6���bݙ����3~Xe��|��πn�P���e4M��I����z6.ӣ:C����=��	�m�ʵ�_XM�gL�L~q�.�M!BY��^|�S`��{u��˿�za�8��/cԛ�7�zO��P�{����ϛw-a�gI�M�����s#Zz�;�^��c�poh��Ф�wy�(��p%�^�y���2��۞���G2�YJ���)���Z�����S%������c�h���ML$�e����܄�Q����Zc�)�y�oJwb&�O{��g�C5����������v/=���8��Ov�5w_e\�jX��m�2>ܗK�hO@�ja2��3��r>kam��D�j9�f����^7wv�Q+����'����ү���p��p�܇��a��)X��<~�o:��K�cq���܏���m����|C�V�H,L��}�xmE@�ZW���p�����P|�㴥��3l"-��G��eg��6��L��ar��T,5����1�2�RZ�N�$Nb�l�� ]Σ��r(jL�$5�~&���;us�[�FY{���?���2�dh��T��5��,���~_��r7�n�����gH���K�Կ�I�͜��V�`���Ȱz��/���b�Tʙa=KK^]�]�������ZƬ���� �_�{P��/(�MY��b�Ic�A�5�~2� ��L��쇚�0�MQ����U��|�f�yAX�O=��쏬�a>;�b(�{pD��8F���6���i�/CP���E�z>��6��g礳LY�-V�_2>s��%Y�眠�4u�!�S�}n;u����swg�n�~8J�o�L�H2�|T9��K�Y�Y��@��R�ޱ0����~�p�r�{�z�H`�!����0�<��Tf-�Dǃ1���<$-<GT2&�Z��� �c�Tb�8�2�P��Dvb�̛r&��U�u�A��&q@n@Ĵo�2�O,lG�2���Q?��h$�8b^�O���D�� ��`a���X3{���P��!	��˰7ϰ���h�9�vyJ��%o����01.�/[4��9�۩�����h�[��_<�5^a�%ǟ�,\���o��&��Ȗ�L��Rw�z�?�cd]�p���1A��G��#�ڀ�RvN�����J0���Km�S�K��c#���{���vD�;U^��C�T7�R�&��UG;c(�t䜙��D����9RO-���e�� `�}�m����2����9�x-;!����|<ؤh漷��iq���,m�g����&��E7>���,у�&'09��
et�e��HG@�N�$i�UGM�Gb�+��n�?0��B�b|�h�ŕKG�#�*`�����
��/"�A�N����o?h0�3yiA�t��s�� Y��bħ��6���rE��޳���JOÜt���� Ҥ��̑�^�P� ���K�S>g,}f|Ǵ}�ݧ�MS�ҞaQ��=�L�G�YX�̯O�i������_��Y�ɯ�_���;ޙY/��˳	Θ@�J[^�P+7[1Z�T����wt�Hi���}��ke�";!�C:lC9�jST:Y׋M�o��Fnn?�?��}�9Q����;Ot�(�����d���u��NOq.#+M��� ��m%(9& <��óZ��/H���ȟW ���:��0������׬3���h�������(� ���_��&��t�M'��ݨ��"|�HY�O�`�٩�mS	�o�pv̧� ě����t�#��]���
���Ղ��&{�3��\�DFn�d��_���k�|��XO���,��<)�N�u���e�p��[ez
�1ü�a�xP�X�:���-�m)�3���8Kq��0x�:����}}SΆ�(���΅K��V����_�(�s@�Q���΁wh��&�ޖf��?���*38��?�GA��u�F6;���ӯ�[��l9�d�����������uC�~�t���A:x]��X���oJ�m���EmQT�Ħ1����gd�K���ir�t��3EW-f�q��3^	=ܫ�t"Z��*�F����ubS�1kj���4�bд8w@�D��Ñ�g1�[1�Ⱦ�� {�{P
�x��j�����:^��Z��-�$���#6%ƭfpH�M��$��=�ޜB����5@���7��]Th���$���ܿ(S����B�ؽ%;�� y��U��6�2�O��W�߻q���</��	1�dAP��H�f�R�18��]�F� cv�H�r�|�ͬg��4�s� ���8���G�Yevgt~#C��E6~}!��f�����ZXQ�šc� }Ȯ�����߶�ԣ��w`���<�d��#��x��,�N/0/�����P�;��@��?λi��E���\��5�`3�������YQ�c�j�#��.�7'�Fi�F8�Z%8X�"B��<�ª]X�z�^�|��y����êk."1�����TN<u����[~e[���^���PU���!%��pW���@���To�B�{���С�L���
��!Q�n��2�<�e�P��kf'��V1ֿ�͜�*z�Z;���b�|��\�o��-���q�7��V��AE�����;ّxپ`C��NoV��F�x#�wN�K�.�Rt�����Ƣ����Z��.h����o5�y7U�/
���v�uo���9}=q���Pͳ�;သ
�T8F<��,�2;�}��?{�ιǐ&E��b��4	\���C�@Hw  *��h����h���/����(��\t��u�}Q�H���`sm*��N�7pM��Q_�w^�����Q<\hV�H	y~B�F'f!�J�$���G�%���)=�y�LT&�V2, 8��3!�V�Z���2����T"k�gNy���m�+{��D����ҒK��2��f�]n쬪^����aoPʤ2�_�_r.�`O�&	�VZz	@�e��_�{�Q�l>kq3N��j��d�C�꿽>���E�z��q�&C�P�u�����X}�jK�wm!6"��>�m��"펳4�gC�b��q����,w��ڿw�X��I��M��a����+j��s�� ��I�b����ޫ]���MG����C0˘�����R�7FP��}d'&�y��ƭ-�o·a�GF͙٣�ׅ%���ԝC��l�BROr�e[�-����bl��v�P��؉e�A�Q�feǍ��X���:���\_��F��{�\X1��_%�s_�|�8Vp/�a�ͻ�F�I�6;.hRa0�� ��%`����E8b?qr�俒��4!�\*)u3;1ߪ��H��Ic��4D !�^�^Y,���r�k&�4V��Īva���mݱ�f��*_�rn��"�H�61�+�MwG$cW����cY]�t�����h�q~b�A@�wM�~�Dl۷�� �b#%���!�Ѵf���_��� �-��l|��Z���QV����"��������1Kyې��G��#�״��}���A����/�/�޺�kV^�_u�������Yi�B<v�箈�h�xбP��:&3l˫�pv>06��1��y<�ɚ���-�P�>��j(�QB�j�o����h���/�?B�n�a@��O��g��ǜ�w߀��M� �OMԾ�sW��r�k8���*��l�oG������)G\�5�;PA>���?�m;oI^�swJy�@���b�y�?'�!�!, ̭{��T��}w�~w��^h J�=�kU�__���s�t���U3+
�)p�E�ذL�zr��O!­��cZ4O��o�2�;��)"��A�t�yUO�����8�m��ӦkJ�9�J�m��t�W)m�Q �tnχEߣ����Q�Z��o�s&�c�b�_'+�Z�����D;��za�fy�+2�طk��2���r���qY�TKd�j$�5
9D��Z��������\]4��7W%5=6pՋ��VY	�]�ŀ,���L��)��؄u�T�����I�6Ϥ�v)+�T�����Y,V*7N�S�On���R�$���t�3 b�h�?�O�nu\QD{R��YT�N�l9G�Ќ\;��G�}N�ؼ��u�V��"���Lx��~O	q�12I�}z�yL�RW�dy��Z�\�K�%�-FF�`� G,$�Ɍ>Q>��U��]nU�����p�ڷ�[��$&:�
�WB�^"C�JosJ�a`���#@���%0mٞN�ָJp�#ŴK�!IRG?������dwW�:���v�O���ebu��w�B���;���S� x܂r �_{y[y�RLS}Y�[`3��e_�lC[(u�Z��0��FW��ɿ����� ��f0�ZТ���!1ƣ[��O4.�$�`��E�t M�6d	u�{,k۱��
6���YΧ�x�r}T����YX���}q�(����\�Fa��?30;��윬�/Bj�uVK�b�t����(�`04��o��=�hS9�d~��;�}V�i��q��_e+=��d������eTS���JI���Gb��2��v��K�O,0К	;	'�2?���-�4�m�+C�$�Uﴺ�h���
V�$���ew2K�l��G"���}��ߏ�g�cQ�g��a�
�^�c�nb1?ԫ�v����V5MԆ�Q�$9;�����	z�ٸ��E�s<����3�2)5�H����1萃�L��7L���<p�R	7�[��'����mH���5����xT�͍VK�Yj����M{vu�Mi��H�Xy�O�8�P��'�	ӕ\��*&ʡ0��*�~����FB�P�qJ������G�V<H}���^���g�7AFY������i��-�s��<�0[����>��|��Ȯ���F���^�*�h"wu�,���ȣ��-`*b�}e�:EF���FC������q'H�0}D`�Q�g����0g���n��ou}�Һ%���P�}?^����u�\1���kr������\e�LQQ���	��T�*\:ę�y�܊����G�D�b.���ce�g�	��p/���Cc���D2ε�r�����f�r�8���(�M4	oՐ��G�<{��VȩY�(Ȫ�ȉ^���	�{��UMs]����:��)�~�K��o�ɶWZ��ô�M·� ���Yiܕ቞/�3U'��d��A��1��M᡼��;՝T�n�+p�-=�pj�r3� �5c�d��D������!(�
�"3/�^)u�*�y�Ӫ�����j�!�����FbFBi)��A@Fʢb���\�_S��0h%Ug՟$�>�4i�Q�����+��L�nS���
{�*�2�2�o��4���s�=���`���3��Y����f�
5Q�i�Ĝ�1�:S����ܜ �Mwh'�`����.���ݘ�o�}q�� RN�|���&Hl�Z%1k��q26��7���a�����?r^�c�U�j��i�D�:��I�X�H!@0ۀ:)��,r6����"頷�jA3��\�C�ݲrnmN�Qc|���㾉o�4�(	:� ��Lgxi���r[�&� ��P#�a����rfT�ܠ�o�y|B�/�ᯏ0U��>�=S��������T/7�L>}��-d����V��^�y +��=j;ꐩz&/�1��,�;S��d�X�4ڮ��zA�.ד��!fI�!6f�q��F�xf�(FaS���Z�a@ �]����ݸ[�~�uX4+��7���4��{z�t_c�ľ����	���5|��R�=Z]|  Y��yD�TA���iT�4�<ڽ���w�_�s	V��s7�Rο�Hjg�#�60��¼�y�n����������42d�JZ��JZI/#�]�ng���?W�E��KkϮ�]��+�l�=�UoҚLo���}1��8�V<�=GE��^����6����1�J<�������46�[�a����r8q�������������ko����o%��ȋ���l��P7��y������c�>b��6f�� ]�	��7#��%{���#��Nn�1�{Li�#�/���<��&����#��&�_@�� Rޖ:��LB��}9�m(�7M~`/TO4"{w��9+l�9�(7R���z���G'�Ż�B��0�\b���d�U O��~X|�Z���w�1|���]����PX�[���
PS`��F�M-�ܚ�v!�C�_%.���5j�I����N��b͂�K�*�94$f@J�J�C��2o8���G�Q�
6��'�����򯪗PIZ����oQ	/+a��}h;��S���s���"~#�]���*����?�S}D>�7�P��bV=>P�_ϗ� �p�k�+�عV/ƊDkQ��)�$_"	���s_AO�n���n
g\��Q��tv"� ���1��\�+6萫�%�i�fI̳->:.�(��]�z�s�:cHLp�ʶ��q����N��S�4U.�uy����Ac�&jO����(�bk��[ARSk��h&y��:���B$:�S�S���W��X)x��gd<�����Ū�!x_aSI����l���<#�Z�A�شhη`�����H�`�+�U4��]������x"����&��P{3c��3�ϧb�?��O
&���櫏Ne�>��ã�2`�I�䒣�E��r����]�:�������
1�����x#����u?��?����O��#0S��@Tj׸.V\��$"*Г�Yd"H����H��,{���5m��N�#�g�5c&#��L'i����oٖ`��~��X�P����\B1���B�RT'��'YPVqV���\�W�P뙎೓�2Xp�_�yJvQ>ݽ���A���#�u<�v�dwMw�麮�4��dq	��<",�5b`����ԧ��x!Ճ���s�*y���i*~�L@��(Z��A-FȄ�Q���������2�*��t׈؛��t�Bn�sLvV����T8-��H�{������Ð aLY\w���e��G�`��A����k��讌�
�5�h��2�od��B�_7�pP�3�Ӳ6s=�A�m�+����,�����e�C,?`�*�1�)�xV;�"}E����W��1$J�HI6�v���o4ZWi��x~ou��A� *����Uҡ�?o���_��e�'�+���eTQ���m-���zUf"�<B�5�����?���}�MO��~��t	��N����O�;���2���'Bw��$тR�v�ńˉ}~#�۱�*GDb-��25tC��sx���1UtrѓJ�1H�|�\\'��E���Z�5��w���F��S����d��̓Q�BnPk���󙩉k�� =e�1+�G�拾G �����j���j�F�P��jt��V��;=.���x�=�ދ4�*|�ȿ���c�;Ir�S�p���*�����;5�GS��bYp  l!\�R��t��^ ��������;�{��>�|۾��0���wR'`�g��SU�ˑ��\[��Z���ra�q�n`vL� ��g�^eK�0����U!��O�naІ[�0���� ��\�3�l������a�C�r(aOqf����۸�~��ܦixKo~��+I��k�!Ӧ�=���#÷�n�%�+��G�VU���DLAep�ɚu�p+�0RfU��(L�_K��,�����{�Q⑸F�I�I�6g����LX�m��A����$As�m_>�רT��@�"��ԟu��!�\z58H��c)��U}�ٯ��~3�(�c�(mX|���s���U�g�@�PQ}�?�}۱�F�d"��Z7���#��8��V+L
kZ�SJ��p�����a�bW���\��,ya�U(�+�ԍ����<������"ؾ�6�ѓ8��j"��Q�|����7]Q�����@q��~t�u�pS݄����?�_ÿ��L�v�lc��Ԩ�T8'G~����*^x��9�7At�5�y޸���>0�Ŏi �Y��q�pYX`�;�Ɔ�;ypĦ��鍞�}N�gHE�%����?LO����3(�~`��}_[�ē�P��;�N5C;c&��=o���p�����~̑Q��S��Rp�������Z��Bj���H�[�4�0j$��,� ����!��s���3���7�$��|���2f
��T�4N�8i�Z/�u�f@�k�u��.!�e[�Y�������4���`j[=����Y���~	�o�(��L�
b��a�ҦÄ�+�B�ETt�_&j�k頮�y���Y73+��}�ʊ8��ڲrT���"V�@�rK<���ݮC$�w��e�:������"L�H�4!��м����F�_�U�j���g/�72�}���k��`˿�N8�Z����3Ү�'�1���W�:,
�x�������0KAѝ9�[��ڊ�57��:�S�f3��M��RTɏ6�������*P��(�a�����񼊈��]�A1�B�ߪ��P���9�����W�A��X�����b�3��+�pp`V���7FL�RۅCX�T���lV1��Q��?�+��;��N!�PW0���r_�[��S_y}�)�|tm�Dp�8I��dj�s;g��_IZ������1~ǔC��q9�S��p/�X��a���!�j����m�#��3����Zp5���q� ���ޣ����ݎz/t��YgL&��C)SÜ�֑2]��Ю�Ǵt��);*��q�!�7�[b�^�ei�/�	����E3#`% K�>�>�&�LBE:|���i%;ݣ���O��a��E�yEw�O����ї���� ��ݍ,��Z�<(����)W5�� i�xy�!������zW�,��5/��>B1��hԪ��Ո�b"�
pd���t[���j
Y0���svD�e]�Ӻ������գdPEoVGQڮz���_A��X��D"?Ƃto��[E �ʂ���d�#�?Z��}`b~�"kZ]�Gotf�mx�Q4��� �%硃��	6lG��E�<�H.�_�!9�Ͻ�uu�r����x�C�)O`?�ݛoI'|�q��/9ᰫ3S��3}�2h���b����"��v�,������w���Ď���7�<�.��bԲ`�� V9?������n9{�w;9T��r˙5�1�;+�E�9b2�g�빛��5�+Ͷ�R�WݷS���#l�:�z��oMZ�ZǛ!���G�xZ�?G9���^����֛ivWi��e�1�����/ep�g^��<.�`#���Ɓ� �_�#�s�S$\.Z��l�����fXL�B���DȈ��v���ͻPjȼ�wanyؑ�Oz���8��\L+�:�-n�-sW�W�������h����[4PV#��jDpM�(>�mɴI-Ũ���-��Q=�����e�#�M�dõ1��:Z�l{ǿ_[T�s^{yy6�qBH�]z<%���Y��h�����N�0���^xyh�������_�k��~��� ���bK�<v�$*P��{�=���p7K�G5z=XM;���<�f���>8���$�fFO�����7PQ�Z��?�=_u^�Wn�I98D���������ij	����J4 �C	+�j�4�|�>rFC~�7�I�l�ʼZ�*�~C���d.��<�k'Q�b9�Nj56r׳�OI�'^`qv�xN�N�h�U\\���8�^*��ҫ�oi7"������'Ү޵���W���Ϙi"��ہ%Vq�X��@�K������O�O16�%�.�m��5'�� ���j�`�.���� �)�3X"�}��c�s*��*�v/��L�©W���5����-�Y.fM�q�~H�����S�'����"��ď��ɲͰ c2�+EOǕ���P�lf��}Ƭv�b���TTP9���@���+���w+z��Y����e�)\�հ��UUd6
���1>�u!�W7�� �=R:��ƏF/ V�d��Rz��J�9G&@k�^��\0�!q��hf��~,I���ؘ����S��(�-��9�bd���yO��q%��;	F��P�?X���rץ����h���)�&�{ �{Ե�f6
c�����z�|��;���B�v�.*A/:�ж2��&�j�e�;[�~D�g���@��Ä溅��?DyD�����1�2�f�پ�R	�'��6s���l� �R>�g5s��iX��D�	��Unm�
'5���O��K8|%x�c���a���]KA�D��k\pګ�mv����d�5c�b�
��kO�^�P�����99S�]w��S7?���K2���2�@8)�M>��u��z�m���w2��Z��d�v���d�s�	?4�����o[��R-]�d��� ��B,����h��K`�&��d_*X"�i<�H������&5^-�ѴQ�ZI��{�n1�7�	��	�J�C d�9���R�E�;G�Q/�8$~�����&t.������d�|��ˣ����un�	�'�94�Wj7��ݾ�O4ǧ;�-�2�z��6h������Ͷ����Ib(5�e	�S�K��cW�fP������=���v���	����Shz�b��(�1�W�Jc���bA���A�gK��Av��"`� 	��P?N`,���MF�/Z�6{0���g��9h�0W�Co�Ah�	"���fAR�'(;(Е�W�����>��/p��j�lcL���Q�O�cWL��*Q�W5jmoIg`<j��?�$�� ��;$�ϢG�!P�ܦ��0G��	����<Ѳ=�JXN4�B�ľ%~��y(�!?�*a7"ԕ0��F�*w�6V]�ddTc^y�#�Ck��u��!���-�,s��,�����4�V�Αe���F�	��R���#����[���ִLJ��t6��E6`��^�u{�w�2�&;���e�Joݔ�uc⣢�ؐ���F0ۯOe_8eB��L������Uk5�E,�W�����q�R[���B/:���ݗ��ş7=��	H=U��eL�l�H}H�]N
�����Q*?�������P/��?�E&�Bo=�[�;�4 ��3�-�".�&�R�[r.ްIu�ﴏ��D�o.�1^�E߱N[d�h1/�5d��j�A@9L�?ͷ/���7 L��� ���t��@H�I�̇��T�%�(�__������+[�&Cd� �X��j�c��C�z0�
c����ze b�sy�&@IHb�0�����b�$�<����L�ޝ l�\�Ʀ-�9����`��,�u���	�[4����נ���T���ź�`{E��+8nҠP
��d�'F�=BYx8�yj�y�Ǽ��C����TNe	)o�;M�cꎯvE�d�Ҝb���/�
� �G�m�̯�{����t�V�h&H\5Z.�p�~:*���F�� ̻�q�D)�Ѫ�f�JE39�aa�u��<S{M�Wt� ���7F��Y�ik��v3��a�`�Mbd��B{wݗ
׵�
��l��Ɖ\����'���f�6��g	N5�p�V339<Q�o�q�	;q%�|���I.�8tRC3��U�F��4�h���%G<�M8="u�:?�;�F���m�;�������LW�}Ӂa�JM�g�Q���U��̀j>M�iVe4Ǭ��1��
���ɰ�u�p=D�'���\���T�&>�O�����}q��J�'�V��
��m�S�0q��y��+���� ����դ��;��fF!�^,I����	����R�;�Hv\��/�$r�������)���R��Y�p-k���7���2Ű��e�(�p��9Z�e9#�m�&��ͷ�E�����^r���9�y8�_��c-��$]�Tj��@+�	���|��`
Ѓ����F���I�Wy��Y�V1�5�kl�}<����Wv
�	��9ǪGQ���^ws�\�N.�{���'�̰B�� :�~P�
*uq��+������vqV��������+����(�$��X�n�!4Uk�F-��/��'�ԕ6~�m��p�}�w}�~n,$<N�=E����-g�ØCH:��H�8Ax�̡�I�ݒ=ϐ�I�#�@R9:S��4�T�j���1
���Z���ס���fhi�^��+̊E���G,ggu�}U��m�"4�'P�^;C�ޛ�w��\�dH�O������n5��֦� ����8��Uܝ[`H�Q����e"�j1�9j�*���/���E���ȨH���q�x����n��? i��#]�9:��ř�O�g���ljz8������N���"��.����1��ZwcT���B~�юP�/�|&��s�#�ԞpG?�	�)�&�ј0�qf� !���!��L�(��$�a�]�QO�N�9^���Be�v9�L}���-���!7sT���c��)i������D�	m��Wq���Y�2�8mb��W�o�z��Z�O�n_�����N��ƀ���ky�	v�죅�^~d��M;y%����_6jw?ۜE�^m��=>֝����略Si����}n?5�`DU�!�O���mo�t��n����/�"8�k������v��!���]�P�.x��y�#�bĒƣT�"��Nᮂ�ά�ƞ�Sn8C�TT#�0�t}HS}� ,	�m{�#�X��.��7�����h��m����0��m g�\�5u.��6�y�����n7�Xsny�mt���a�X{��i`1�}ܲ����v2�)פߟE��g���1~ӎ�ϵ�!��|ԃ����+`'������MY��3�!�n�&c���@3���D��K���Β���Z٪Xjr����3A% �@��UWi�����Q|hr�7�C󁪊�/�3����i��6W"�uJ�t'q�b߬C�D0�x�F��v�H ��
����n����Qyl)��8r�����s��3#��zq2x��i�CיW�A)P�@r�|�!>�|�_Q��������ˤ�w�
�lP"��3��s�$��)	o�s禂pn��gr�0�TiU�:�{عc�I�R��j�����%�R>��vy�`�+��$�j�M������:>{�k�1O¬$�%�{ʡ���Ne�ھ,�\�IXu50����F�ۑ�@��cd�����:���U&�K�W ��b�(�Udx��p�q�L�6�m�e��>�8۵s[(gY&X�<yp5��>�Q3U����uh�G̾����T�q���G�� ���l��#�J��J�t�x�3�{�3l�/[$8+k���77-��6╪�Bp�MN�3ʐ.{2uz�ߌ��?����cY�_�vp��~phz��)��b��8�H@`� ~U`��9R�
D���� ��L~P'1$����`�q�F�_��/N���Nb�0��g/����T��X�a�%�g]���P5��s#�U�>��9 {.�Zf�F*����Pz{��h&/�`��dN�5�H8+ E3��e)<l$w��Ũ��&��=���b�+S��d<Qk�R+��M,2}�nC�	�nyy��b�GD?7���j�Iz�=v�H�Ll[�xK���= �a�f��t���k(���UG�xU�Q��1�<��ɋ�)�����.������R�>�g��Vj?�l��%��JU��6I�/r��R+3��e�Z	(�>f�>�8h��H�Ej�q�+�5<�x�+�IG�	�aDZ<���z�����B�g��s��	��b!�{������"��>}$��w������Ǔ�]$b�E��3�=6��L1�R/����m#�1nF�72��*�ZR�ygO�q��Tt�=c-u�x݌�p.�}���8�� D�`3�������q�%ך�,�ԓ�jN�Tl�����c�vc���
n��t
�x1Ѽ�5}���(D=;�CP4u2�W%������y���7ٰ��	�T�m��1.5d���b!��{*�+����mB�)�t���.�`���Ww�.���zpU�90��ݔ��}�%O%y��Ϻ�Ng_Roux��p2��3�,�rR$wj����W��i�}8���}�/:��,�5�^OY�_웖��DANS3�Kc֯ 1)4����_Pʤ��zd��t��{�f���o�
��yq (N~�}�Ξ&��_�~�;H�	����m��Ϡ?.�٬8Xܟ����=Ws�t����p.m���@w����U�"���m	3:5�$&�������C%[I���h�S�S��c���C�~%��Ss�N%���@y2�pBM����ܓ�hu����&�,�ݜ�'��&�'.��q(�;U��51?�9A���GO�
)�~�(3J�6ab�PC���&q�(7���uv�B���Pe�:��7���ϑ�R5^Yf�!�L�%�q�܌���ڤy��j6�%�/y/A_���J&��{_��?�V�|�OdU:pq�0��Lmwd>	����E1�������A+�&�W�g���X�"�,�{È�����'�V=$l�y���ЙV�v�Be�)�8*���@��u�����ar/��yP�CS�f�׬��nb�OY�{�K��ب����#x6Hw5���m1R�yZ̈́����p�ERx�u'���0Vkw$+u�[Ta�������۰��kk�N�7�ε��l�Ru:��D�WL��nH^S��g׭*3���y��fR��N�Uo��`�Y(ڣL�� R�q2���/Z^��b\�L���&�HR 6I:F�w,�ŋ��ؓg�X�V0�4kMP"Aa-�lF	������U�[�o��I��N���TBj���\��x4!���6�esS�U�DoO�'�}�a��k�j�_�$�L���O�9��dPݽ��|�@�it���n#�M:��_AI���^7����p�v��^��� �H� '��
�X�$PN��Un�`�䇡.B�;k�V��[)�9^�f���۪�N9���ûdk :efD��y;����_3�n��p���� �8�b��Mu�ё[�XQ>W划���v%SQ���c���h�`�����Q�ǈ�9~����/������l��&�U����1,3�|j��X�֩r��}�K��ʐh6z��;��EM�W��<"��{����W�g�·r�K��ٌz��,`�c�~�dPr�St�B�ҬPNA9 ���K1��f�yW����u�a�xC���Xlɟ��]�Ѫ�3]���ޑ,���CP?N*[v{�e�nA��C�Iǒ�0��!2p�H�oj7��{"xc�g�X�����G}�.ޮ��{]���O��6�a���*�Q�q�,��xp���*��`���v4]�	n��|9�o��񥹻@�Ͻ�i%X������WB�Jy��5_��L>a��8W�Ʒu(�FI�|��<m(�1��`�Wf~C8^���R�S;O�ax����s��V�
�� 2M��؆����yۡ-`Ŷ�㫳�0���u��QD�����[y'��Ҫ�������K{qC��+��_�1Ż����Pi+����ϣXH��ٓ�{D!�4��L�K��`¯�b�A�j�����ل�+�'����0.��L�?�sV j+�\[�År�3w4TSyiz��*7�k����?�>p`��1bծ[Ք7]5z$�z��^ch}�~�&g��=}��ҩ��Q�E��/��޷l�_h�U�57���T�q����O��*��۪S�Y-�c+�\��;IՊ}����t��lЄ�S�֠*ȍ����+�z�ޅ�E�o\�	h��з�ifLo�A�;;�H5�#�G���TvmS�)\�i���!3�- !��x�P�Hj��i^���y�s/�R�j���1�0���Eԩ�"��j�������9���^'��d�Y�t�����~7,m3�]�Tw?����H?�Īuޟ$Ŏ}f�W�2uX3�*�� 
�qڮxf��>A�����/�	O䈹hvǉ/�G�bJ�L�W�9wi:0�S�f�S}�����]��w��v��N��]`�8Q�	���\]z�q�������YJΪ�C�k�ɺ.D8,��9��g����|U�A4s���h@�B@X��5 �rm%G�R2�;!9��Ī ��r"wK��:���P����o:L��R�KB�z1Ғu��)kX���0�p�!ٔO���h�V�_x+5�&h�V��G}����X�>���=e���,cz\	�����2""Ep�W�-�!�w�ǣF���g-�
%��dhi\~��ֹUA��Or(+ҿQ�����C��{m.�͵X��������0��V	��	%i�"+���T��[�a�u��)C���*%g�n���Э�@	Z��4����~5I�$�w݁	u�O�-o�#��cE��x�����7c��C��i�Z�6B�n�Dd�!�n}�z�~���0��ԛ�#�-�!p~�GH��vo||?x �?Pਔ���n��?�8�<��[���-��4��<��F9�n
�e���M$h��c�k��1H�����w~���T�kj5�S�� K}��O?�/�*�5��l-=�Z�6:��Q'��������z�{P��`lm����\�.��Л��u�s�=.$:)�3����bpI�z�.k;�7i4�ԙ�G$Ap`���d��%�M�
d��D"�[��b�L�e��wo��1�Xo�+��T�7�q���N��@�U�q�)�*��������%��S���
{�Qr�JL�NE"�Y�PG_�gk�Kէ�֗}!n &z��+�tl�J�	bκ9hB({T��*��p�5q9�衢�;�;��M,.�MwT�^5��%~^��'ҡ9�ķ��$���Ħ�Q'�ۆ��Jc���^�����Μ�l��������#�`����G�P�$�諭=�>zbFF����b) �R�*Ej�O��3�?e�fy_���N�t��X{�]���x<Q��a1��%�Uͽ��F@��}\j:�o����ô�(����+��;ܴ��h1i�o2l�"��oa���
�b o�Na�/�;���<�̚I�믌��� ��Q۰�}����"锳�Y���n:�T�?�CMW�6dO��<:?��I�i-���v�Eu��H��f�������u �)~�Y�7'@CSTu���Ϭ�=�V�� �T����0u���}�#��	*��P�����	٪�S��ǔ�_6�@Ԙ��-��	����0�x~>��A9NKt٬LPb*��3�vnM���͸�+����8~�^˹��b~GU+��װϞ��!��׸�[ԧ�o�Y�Z�bW��9��g��λ����፪7_�ih�X��g�E�"���0��X�fk	����o`Ђ}�Z@��9-�����iX��%�gg}q�F�~	��e�����6�VA�+З�����n��^���zͩzѺo�,Rv�xD���
ozO��`޾�B��.�3]I5ю~��Ct�S�.Mr-�W$nOQ�/E�L�F6��8jz��8�l�?Z��l����1�'c���(�������kpE;Uf�벅徺�f��V�2t���ÔW�5d-M�Q���Q�q��� �iWT����5[?L�Yq�q�/j /��`�����$�ya��ΰ���$	&�0-`���(�q��̻`���n�I�Ɯ�v=[��mn�`�o'��	��;EQ,���&j�7�X���o�`�R�����Y@Pb�	rj��_�wb���� ���N���v
�aM�3�L���?�x.Ă�1u��2��(, �SM��`�k3�|��ݑ0��IS��Ò[��b��r�"��v�a��dg#f٭��-��v�}�P�~H�H�36Hmȳ��=:���N��W713]�"�ް
Y�W�?��q��X�	N}����B�)�>~R�g+�#̚ʸ��7��3��J�aȓ�`��0����ӽ��o"5$��d4̓���`)9�ݛY:@D ҍT
��q©��s dЮ'�~��Q-�?̅��DA׷j�8�����<��p}ӝ�ݬR�i���M.&@sK��Β�`K%�G��T����!?�Ңq�b�ʵ;����m)t�xZ�ZI��o@�B�^�$���>Q��7�_��i=%h�S�����
�u,�9�|�$��PY�	��=D��ȘŊN��B��D�҈Ԓ<�WO4���B��辸\#Ǡ���Xx���<���T"�3l��`@�'n��Z'l`���c�ӌ��a���(*=��o舆Vrm`��nX8SA��KX�bkv8M-� ���3鎩���k��Q+;��c�%2�:=[JtF�4�����6�s��bP��;m�(���["�bd*��;��L���w��w���>w���8�e[^=9L-<I�cOV	�v�NX$Oq�Pn��-�V˽��(J'�l��b�D`0­��<]���Tu1%
����0߈q�C�1�]gT7@��Iql}�y���9�8�i��m�=�)TL�uMcFz�gZ��f��2)�����l]{"�i���K�2�<��3K-3�p�N�}�r~�l͵���SJi�FGt��7%ޤ�0�]H��ﶊE���,?"���8h��q�f�Q���"��z��Wz����(12=�*'���S^�`�z�}��7.(Ae	*t���	����@�%��L�w���A�ܰ�+�"����^c7j����d��P����7��!X��2z㓅��m��+��9A1@�[#�xlf^�c0�MX��g�]�K�0���\�z�`#�y��ʿ}���)��HC�N�wP��@׃p��&�MN-N�U:=X���*I��˯���U�u��N\k�%"��k�R�:Ye�fj��j�ܯ펢����� ���X`���qc{^$RL�'".��t���e�+^8����Pnq�Hw����Q�����	ŽW���z���,1/�Y�׆����ݖy�\P��Ā������W�4��h� \]m�y3Y��Kn�3<@~��͂j,?����š���6_�T��V�t!�P���iy��-��A�l��W��Y�6�.ﱘ����]�4/��Y�i�j�l��s #;��f���?s���5����i�
�`��V�c��+�k�W��ⴓn=��/\�P�+̃Ao"EeX2�M�`qYtX�!H�}3��w"��5P��f���ak��,��I����ޓ,�Wi�?[P��î|(m/yJ2��~1E�\��Ks{)>������H֡��u0��=����U��{Z��.~'{, �$_�PY��㎥�?^�K��B�z+Ncp�+�m�_�(T�Q����%�2l���%�鯸�N��%�1�e3�@kd{�SH��e�jy��Y����k"�(��$?D�ʦOJJҎx``�8��L��m���i�p�ڿ;��\WQ��h<��PQ���@�z�p��;�_�8V=�,p��xf�{�@C%�[��j��A�� �d�T��X�_��d8^���hA|6�P���a�a?�h:��W�5�RlR���ObySQ>���b������Q������TA%��r�����I�Լ�+����l��w���*�rN�sV��������o����q��k#�]�w��*;��f2��	t��h�N���eo����v�q@:�$P΃k�[�j�m(�Q� ����8�/h�p�tn�����:
���^�H�q}���־�6���@'|�SU'O Z�$�[Ѽ��F�W�R�(-|����\L.Y5l�eg��&}�)�����-��_7E��n�rj|���}�_YK�ھH�`D@R}<�R֒��L�� �� �>V���0'��� �~=f�Ƨޠ�Y�Ct�sv��r$�rZR�7��7���e��{TTV��b�+���m5Ƃ"gxLG%�s$��X�~ ��V#���A�A5IZO�Kq�bX2�ū�e�)����頨8=�R�]gJ��J�r�f�6��6H���;��>!3�����!��F�m�zC���	XN����Z�t/��[�KQ��uNj���	H��j�
Hwk,�Q$e�4/D��n�/�<e-h^��������$�w�<��x	"�H�kX�����n؊n5���YH���h@U�Z�A3S��z.6>���7��@-
�Q�r
s�<��B�3YW���
�x�p�=8���(�y/�D<���Q�h%����
���$<����,�d���v+���#SȮ�����+�̂��΢ʤ��c4�#䨌K
8e��]�;�%|e��~3��vp� /��gS�wI���o��z�?��bHj�S闯w����G�D����	��ԋ�xk<Xli��G��<�O�\�$�����B�3�Q� C�B���-��f/�ޙ��&�qB��$�cm��@@t�N�,¯�����)~=�ѵ2�5���͘��%��}jչ��e��Lh���*[��cM� ��/H,�[���?����k��l�GU ���P.�*�X�ž+%�?�,)��b�I��@�=�pZ\������Vҋ{���]i�~�Qs�Q=�KR��f��Y�]VD�]�§�+�z�.�K(�ױ���኏�o�;B����~Hb8[��7(<���&�w�)\���g(��Y)��JNJ&��U$��Fp��g  �x�T�D�JL��~0�G3�����L�K0��;.�c^(�K�P���I!G5����5�w��H��$zє��� �?V�W�d�K-m-C#M*S��-��nqb�n�r�-w�<�~̚�;ʣ��h!��a^׷�Y��	�F c�Ƚ��� ��e5��$�S�����P{���7�)�g:#7�%�h��w����wN���4�a�1����B{�����>I<R��-_-C�d�ڙį��%�����6����uᴠ���W�K��O�d��~	�Z��c-�-��U��5�A�>�-�{fM�Q�S�`9:��H@��a^�&��4tSҘ�_ܝ�\8|���X\Z�ऺ�A���,����k���ڸJ!�.�-^d�g�qAN�^���5�s��MQ�����"jl���o����t8���vy�9^#\e��N�S�B%QQ��0�nD=y浗�s�����
�4;��f̐�>^�C��q �"^+I	����J��]P�%,t����j�ݒI���!8��Gc��bsHR�J��D�7*w�2�܅�f�8'zk���-0�}��$���y�Ro7j�0 
�Sè����J::4���k��lE$��s�)�a���/�ֽ^'�32q���$�	w$�[��v�6��;�[t�ݣ}5C���M����Ɛ��s2LٺR���n��֧��Ēn!�1�D�	7{/��:@,L���jW]MG���MoY%*C#���-�� 9a���#��-	K/X����4J5�X�����(��[��!�h2g	~�ʉ��D5|��\��L�P��i/9�R���4�,�_����Mrr�݊���FT�`�W�Fk�}���>��;5kC���iQ�0�������2��:+"C[�+yi&	�W�ook���fK�������U�Ş[8;��L�'k���?���A'� ���[j$�J�ڢ9�ܳ1�|m�#^E��҃�2#�I���HZc��0_�*9l�'4�������ϳ�X��/��V}&�ɏ��e�!�-VR���+�~��&�h��ּ�i�i��l�#��ATQG���\{�Q����vK����A�SI�v'T��m�YP1k�n�2`EZ(��>���
w9��j���W�xV��rHi�'� 
���a�Ù,l�W;Un�+�4j�9�ً���ーb9^(
e��%���܏ȔtO3�u��S��E�3>�<j(��I�%�v��O?���dc�V��P�z��u�6��*�#�A"�9'��n��M����n�F�S�B |�>ێ`<����6��`�Y2;�S���4���>�+[���3P-��.�����)�]�b���U��\X+���V�A7�g�ӸUc\3�5���A7��
�t���O���=ri��mӫ&�ˊ\x�L�ͪC97G��#5A�����I�j]R�F��^�����xm@����%t�G���B�wpP$���j��aiC�G��1��Y?�:pB�) {�yA�?vlvpN͎Q��215"9"��L4s��9�f��Y�r,4g	��ؓ�Fס��"x+�(�X�HˆM(d�Ic�\�{�1���
zP�8�l�!~̢��T_8jI���``��d��O>��Dpd�c1���*��/�i���2�s�mv�~w`�;&JOxOT���+ۖ�W_�}��%Y�`
G�#� 5x�y١zk�̕ iokm���mR�O���E+=�4�ԅ�ןb����q��692�B����Uy��!�kX7�d�j^XN�"uj����;MJ��i� �7���^��̤��#a�mE���Ja�%�`���!�->�Gm$y�s)�O�6M6�[��_3�7	���.���t�|,�ϖ����@*���\��M)ܙ�℅�,��O���2�����˚o�������U���*t�b��v���bU�`U�Mȉ��?Y����j�Sbт�=��j�d|h
��k���:�f�Ux�W�qhl��9V�B	���(N=:`/�:Z'�C��0�q��e5��?z�%�(��Q��;�Sg�m�[EE��
�k� W��I��=pD���u*���7��%.�?d�tν�T��F&�	Y����(<�����=���1�ŋ�V�!6	��F�I��n��˰M61P�{��1�4���dB��F/�X�����-Ob��s��y:Z��1zx��>c������h� �ɷ|���*�_s���s�㟬�i�d�F�hԀ��R�ұT��E��8Z=���%p�
�~��S9��=�Ͼ_�� ]R�U+�C�!J�~�y3e/�k�2�`��(�k����^k��E��J"O��>}�5� ����O�w�R^�9Yj�i�5���W�d/�Y=��9
_� #���4W-�w ���Θ6/����&�<Dݒ�6R���n���'�2�{L�B�zj�^{��}�Uo^R�t*X�s����-D�OH���1��x�yZ,ˑ7�H;I|6\��f��oT��\�?vP���������V�z$�x�ZJ��ޱX���^���4�����I�nFZ\G�ZZ��C��v��p��%��\).x7��m\��0������a���L�$�J�#|	YW��7���h6�YN���~��jm,D" �;��,�yp��p`N�u)P$ ��bO���!t�<tYe�W��R�u/C��{���#�36�w�\���n�=^}~���a��rF%�����,�����_��x}��HE����%@w���ӗ�<��l�7\��*�b%H k��BQ�X�&ʤ��<4�%K:���˘���9��f%�<��B�F?�2��I�##�D��a@`�3z=�*��n
\�a9���a�h�h�\ƞ�V2�j�sގл���pZ8�!W�lQ��2� ���Dw��8�9�b�ݩѴ)�!u�ί��������\Ʒ��^�V3L��	�;����]r�-FK��WuA�G����Y���>&���7n�
�*��Db~K�iN|������.�����j?�1>b���aM��TP�y��,Hz�}�U<�L�����#���N���K'��1�o�|�6�[����"��>=R�N��y$2�����x�DS<��qoi�.3=���S�~�
ޗ��^X���rGɿ[�}V�H�7��������b�F{ӣQ�8�Ľ4ĩhٿW���;[���	�fl����>@�U��\�0��hP�vC����;����*�������D�?�6�"UI��0�<��_Q��*A�)�g�Ugl�_�	^M/�/E%�ԗ��e{�<�Q��=A��&��j��F�}*㻆�yh�n�����4�*��.�-���ţ��p��
DD)���Fq�[��I��	�=�"�[�.�%��	rDWy�I	�	K�L��r�*�d
��0���[�3��#:�)&3Kж�Ϫr�0s���X���;_o{�����������ՙNYB߯!�,���$��%3�$��!g���Ǳ|�'Z��� 6�|Ik��̏;HX�(���'�>pI���a)z��1a���x�`7��:��,���$����o��gBU�0"#����?
8���Q\ja�`���N-Q�cB������/�Y1c��YT8ދ Ћ�<N��p�jy}��ZZ��uA�J��<�\|�P+�#7�����Hr�a*]�a֏�tL��$� ���C]S��&��^m���������� .U-h���ԃ.�����y������-�Z?�� ��,*�gfC�z�@V{�)��T+��p�#�~���gg%:�>��"��0�*���b/��8����|ꙃ6�~C@�l`�Q/^㥙���̑�]��#\q��F�h�M{4�y��� N[�!t��	����=h��L�-�*r#H$?�^eԔ 'D��ܯr�w�3� Ç,�| g9�F�ꩳ��TҀ��'�#4ʉ48�����!�����j��.��Y�.✺��!3@���(�<Y�1���Ro]@Mш��c�����[I�9/}�n�����C�)P�`��n ]���n�戬g���SO�����aeҀ�V�~[����ޜ.3���r��Q��
�����<���.�pPT� |k/&@��&���ucP�A�����Y0�������ɪgz����ݤ�%r:�
f��T�bA���������G7~?М���
��V�\�ȥ�x^�a1U����D�UZ�kV����z(~F��F~r�c!������@|�ccӅȶի`=+��������f��"2x��8�mŠ�X榰�������n)TOpCs�#�)�D�uO�\Xzs� �%)������6�r��qG �������D��� ���
��M2b��Q�3+�__&�����Y�Y�T��X�RK�*��ߛF-C5���Y��,�K�Ђ[He��[��?+#�Ԑ���q���i�y�Q�Ω'��c?����ι���sV݇Aˍh�m���a�W�1S~��ylaƄ� :u�I�|ƾ7�c, �"6� d2zWYy�����������(��D��� ��Y���=�9y`�]�wk��N����a#Mڷ���OkR�}�b� W���)��EĖLM��$
�vN�8�{'����7r �+�y�T5�4G�C?�q�h�ӻ���j3%�pd�3����^ff����?n٬��v��KwPʊ'�&��G�$��)�#� �h�'5��g�( 4"�G˩�j����E�=�S�R�Ɵ�����$?�l������u�K�䶲{�\]�,+E:�0�0߶�l>e��}�Gf~@2l�߽�<8k�Ϝ��.�I�sa��g͓!�[�&�Sx��N޸��Œ�@���&��A�#J�g:8�/��0�e�Mm�M�O���dl���S��8��B����0�6B,)U�"W�t��;�VhA7Ak�J��Ӓ /�}/X��Y��6  �v�
�e��P
�i}�ҏI9�D��r�x.:�K�:
B����X�����TR��M���8�  ��`+<�pJ�Q���mn}�q �;{�V�Bf�d�^����^��
�Fd�?���:��- �)X�@�^����>������^o�����^��m��O����0l�Q{-I����v5.�7M	�9����M���U����~)�/�~KҰ�[h��O�@�mɊ*��P6�n#W�2���^l>��jN��ZFP^ 5g��;5�H���%�������bɿ���Ȱ�p���s!ڄ9�|�Sa���~�UL�q�����˽�i�'�r�4�PA����w���w]]��oŜ�;�-����傇��{�f��o��ڂ�x�%"�9 -*�ϣ�����i�ó:�u���QqjOBO�eH���)�C<�ho��{v��jq��@�Y?��@`5:�~�މH���%�Y cD�n#G�f�Z�b���T��ra���N�+�0�'^6��u;V�G�N���^�-7�����b�z[6�[ЧIM�oU0'�XG����e�4��\R�D,�5���)r�N�l�OX��t`���;�+ ���ї�"�:�����x�ډ�C3L`�k��g���BKN�	/�����8f収fu73�K0���
�HY`ն��B���8���]��Z�v�ඞ��5�r����<�'�����hX~.�%�xM�X��,�ix�s�����8�댌��b��v^b�^��+	��F��.�}��Aبv.���Y��g�p�[��D�����ƹN�*d�p�3��^�R�#Kqc�AwլCr7��oX�Nu4$r`���v�_��.7x�����
���xaJY����L��y�:2O���l��͕#<~cY���b��K ��ڊs__�^p�����&��[��n\S�����B�p��7�`(V�;�d���z�h�9ƃiN��0xp���O�����V�b���=8���D\���\A�8�5ԛ+�j�eL�z����oTh�J�]����90��m�E�?Ҙ;~|��΅�\p�ɹ���Lϐ� '��Q�55���u9�D�	��RpQ\���y�#�G�yO�ZoX�c�X�K����kW����|�h�YA���S�]	��w)�B��~Xѱ�Ö������`�L<�P����L��M6g�2�{� JV�hV�$`�f�$@�8��&����X.en�}���vb��Fͽ������{W��-�) �� D����D�&5����s2.�=Hm*��x�'x�������?τ�¿H��n�"D�h�aZeC��,�x֗u�e��M:k��y�h\�/��T�Z3h]��D���fl"�#��l����@�h�C����W�F������9�Կb�UǓ1Ƃ�zɢ�D��D]t��S������o��Y*(e�.�i�D���w��ġǎ�̌i�Z.�/���դE����IV
���-s�1QG!^��m�[��w"u����F�(��������6�?�������C.��${N�&qT�z��2����lt� ��S?�sV����aD��G>�*wS�J�����^~HB��7Z�\vA����g������:&#��QNY�2�iR�M���`r�L1d3�w,��j������x@�E�=.����z?�Y�5�0��6T5t��6S���M G���φ��]�ij�W~9�2CP�Ⱥb@�$y).lG®Xb����g40�/H?��@��C�X J�������ܑ�&�M�*�q�����
�P�M8@�6���]l3����E���{�
\F�ɵ��p�����l�D��R,ܡ\ϵ��,�c����s����1�ut����u�F�A��񀠈Xp��6��<�7��� �������%�3� �Fm_�v���:
&J$�1{�\O窢�;��B������Vp꩛g12��6��Ι����KCޛ�:$?i�;���c�
̴�j���<tj�ZsH��\vY*}���E� B�T�%��������Y����:`w�'���A!!h��QB$f8Ʈء����y4�h�[ᢉb��г�����D�*ʝOq�6�ڦ�z؜k*35�l�/�>ڀ[�ԩ�:!/RqA��>5��W�Ѩ|R�J�&�)ٟ7��ġ�n�M�DZ�s�����*]��0Ԋ�r Ls�P�@��L��C<�#���FtS'�|�W-�q�Y ��iQ
�/�+a�?A׆:�n�"�fN�$��a��4�[;z��ޯέ��j�N��"�9�[�y�E�V��ޗ�� ��v.r_����pm��ȭ�|F�_o�6�Ǒ��#e��0 n">�1���M��|Zo`�˿�W�� g�W��_oϳ����ֺ&:��V7�ݾⴆu\~}�O��t�JY���1�ԣ��3����V��b����+�KUw.�2"g�7�� �,���:�U�h�~�Q�����B�%�A���|:>�Ḑ�h�S+���;;���y�
?����@��� {���;�S�=�@�H��*X��
P�"�JkTv\�Vز{�C��X8�0ʂ�nd��ϭ���شD�ˏ�m��^o]����f�A(���\���ڊ���(��dg����[�6��#����(.I���Q��9;Pwc�Y�W��U~�=2�[�w�v���4�5��z��32���������	�1�?��F<��K9�V�&�I����4*����1$�P��^���ұ��b�S�eT�c��_�W�@�5�h�n�i�~�^4�� ����;��3q��$w`F���r�)�k�(�#s0��r-�qg���"�X+���=��K@��͍��f�C�X��;D
�w�c�F�^xEٺ@Ê.-�~_��a��Xo���)��I�W�gh���/�YPk�,�,S��j����qp)̸����z��!�;�w�0=6��zf�Y���Kh�n�����C�����^���Q�]Fַ��y���yV�ӧG���G�QV�A�GO`�!���dr\��N��|i����S>Z�2B��:�2Uv�+Q3iE5��]D����A�����_% )\�e�����uӜk3u17�
�ţ��.��X���2w����Ƕ�ZM`(%�!�����-+�k3��M1.�����ήVy�,<�O~��+B��[+��'��M��["翧��fT�ǅ����91!J�S&��l}���;�,�* ����%t�t����W� �ѓ#W�(X��5$�d��D;d�n����03��TR#2���hJ@n>�ڻBF�[F�42��ˢ͠\��(�t�i��X�; >?�D�G#�`r�>�a�h�>� z��*�1����(z�5��W	���y4	s?��Qbs�'�V�#��^�(�'v�@���>�M�Q��+��X���b�RgK�ծ�f�b�coo������L[� ��f���˫L�ss�dݏ���������u0i���Ơ�l�ĭ���N���i��C�v(sf]���[=	�=�=� C����J���hl��yS���
�;���2������[�ZO�����}@䜒Bᜑ�c!��;�-��د��J���6��R^H���|YM��e���K�&�Ӻ���(}!�ӟu��V@�'����U?�N��<�
zv2����(�'����v͜-��'�b|WqC�d�璆���.a�+�>��0�ߎs|��[e�f��`�����Fn�\����F��O~i�<��(�H��3p���ݚK�~Xˉ����J]��l ������"���l��Uy�S ��Ʈ'a4@I?w��j+��Ec���;-HmM�\�H�H��oݡx;�[9A�j�K(U�^�Mo
Q!N�rO �\m'�tx�+�$����V\g��F���]�rg��""; <(�ڑ�讽��h�-u�j�s�Zw��a�˟R�;&f�c�Ӧ ��|�&t?�`v�J�g<���A̳��SD&��W���4�n�m�KC��֝�$������m������P23�iOm�/��M�y��VfM�L%�i�xM���s�ŷ���y���r=b�Zg v��mw!������=!�E�����)N��'=[�`Z!)���oX��o7h�+����w(�U}�:�N�9�##Iܴ�.bͮ���ObY���)��W�+��w�����D�6�r�y��#w�6��$Ck6h�M�.	�+}��|`�֕]�ґ���͏��MO�v��9Fyl��zKmU"ɶ*�tض[I��0J2k�S��$ ���h�Ǵ+��x��։|Ğ�h���zGa��o��n�ue�vJ䝡��L5!���B��4�
��k�U��"���z�� W)��4)�~?�@��g������ph���a� ���%���4�]��pd�z�/�'2 �`����ҥo��܇m'�A�Ƣ3MLD��������U�DA;(//Z�Aӗ�.��4Y����ߖ��k ���c�R�����0��{|F�A���r~���>�)N��%~3�n�=}�b��0���څ$eԪ��͊��0Lq�?�d�������P&��[,H��M�XLI�e�� ����4��G���φ�&���;^�o����p(�_d&�^�5*~?�w���K�X�x<�#~�A�I���	���K<7��� �!G�AA/�Brrv�\����{ Wo!�MN�&HaU�
�H�*�CW�#�т���)��'�#] �5��\���ݘy��֊���[�/���K�k�͙�Є]��G���� ���K��m,}�]�C�<��'�Z����p�Z�د����ZIۺ�Wk��_�� ����I�t|�\�M�s��&�u�ך7ǭ�=h�W���>=Njh��X��m��F�a��fekGR{i�*���!�SS��}ݥ��ǘ�����BH-æo6Î� <�#���*�.�X85�&�o�
��	��X�t*�������V.s��"K����;������a%�N]G�Y;��*�ɾb�H
7��BSD9�Cn��)�V:��g��Ůp���¹�?���MThg�P�.h�d�4����G�6�&Ӻ�x��O%�j�0p���C��1G�zJ,g��4��^R9�����C������d����u,.�e�,���Z�}V�N�J��F����'���5���P���7��a���߫G�H U�_�wh���-W�����#Z1�Ij���]�(p��x���{�Da�#��k��5
���/���/����ʝ_�jA��<ͮ3�I��������ҭ�G�����f�*��s��T7C�<A��w�m���j�j��wA����诐��btS�nϵ�ki- �){ކ�h���&�'z�_�q�i}Ѣ��x8�~�,�2�'��?3�C��-�E���:��ix�x\Λ^X16����d$XArQ�<Ƶ��nI��@6Fo;FW���?�{�4{b����������C�Ɂ.���J�?��ޟ~��S��
��/�����m�������U�7],��KلOw�Rw�>�Q`ƺ����ri�X&(�<���'�6%�	W>��Ѝe�n������G"<� �B�Ͳ�]��Jn���z��_m\H&mZ��o�vqL�l����,ڟ�7�>-��è�PG�aAw�)N�w��1�F���.y�j�sG����n��p؈fc0�kl�!�Q&]�f���E�]�<hhXǺ]"��sͨ�.�(���X4���0�qɟ�������F��"�B���ݭ���+o�e���a�w%cז1�Kp��߱+T��eqը,�7l�z��1ۋ0<׾{8\��}�2�ˤ&B��{��r���T��y�\���������U�f�=$��7��~)q��IH&�w�����>��
	k=tE��讪���#�����p*��Dz0܍��i�87�H�$[������ ؽ�8h�P�Y,��jE=�=W��︧��&?0oBQf�،���YL]I#���D���<�9�C��c�s�����Dr�#&럖u��$G|Go�'�&���Hߨ��1P �(�X�*�.���o��>Td����o_�l9�a���m��_�e��XS�{wΛ��LT�;|�✢�o�R�.�����(WmC�iPj�>!f�<����ƌ-x8�z�t]�<�M �®]�Hඛ�lX1�0���?��|��O�g^�L�λ��^_�7"酢t�77!_����J �:.�-0О����[���4���O�~❸g���Im�����1p%��;9A,�,T���Be�M!+[*�w^�g��q�����S��b��n���9o�c<�F�X���K�3��ڪ����ڑ�ӢD�t�?���T�F��V�>=����ݘPr����يN7�ͼ�@�MWhn.�D�4L����$�F#
�fGG3U���6�k�LC���n�-Ym�L��,��h��i�����_ҩ��B�U��ݪ�.����9�f�}#�#y���P�#�P4��6wL9Ų��������e�]�7�,{�suB\ݼ�G�?����ؓ,�k�Xj;B�ռ��@0����������MĐ8"t���G[kؖ�ݙ@#�g���E�r 2qn��`�7��b�S7C��_�v�w̓<�O�f�"�N�X��GW��8��t����Qʚ���w;�K���b��R�`�v�Lw�1�G$ՓU�*�3��� �)�#������Z��&�����!m��R*Z��^����3��ٍ!Ѷ_'NJv��q{�sY�u]�,��[Z
���p@vl��ǟ9�����?v�To(#�z%-�Ǘg<�-Q�c>C�� I�FZ|i���k��R��^i��뻹B|�A�2���!�g_@
	⌖&�d1U9k'`�q��nT;߼�$�D�ޭ���������j�@*,�%V"�O��o��T�4�Oଊf�߃H�_ъ�⁒~z����D�)�p ������ Q\c������Q&�KYW�$ެ�G�(HC��#�~�:,^5P����aҌ���i�~d����2bc-h\�S��.�-M�~�z�ς���x;�5�HY��խ��~:��IB 3,��M�4\���~A�G�q���0�
L!��������-�"S�V���R�!����f��Z��t�a���!R�#�*���.�WN�xr���+m��'C=vl�f�{�������'|�"�H�6O��pN�Jߖ�����K=:1��S2�^���F���ϋ�O$œ1iM���������W���Eo���N;�qQER�s��7? ��j��J�\! wXU2�`}`ip�c�|��P�Se'��V^hjǒa��c(��9H>����OJy?
C����F��|lT���$s��%�:RCYi
�p�Y��1�hn��+m�.��v.zj
�5��N_�^���>�g?��|{tg:/$��{D�����{*�z����m�>d�<C<�=�ޚ��kͽ
ə�����r�Z����N.9��O=���=žX������ڷPp㓿������JE)n�Ծ����K �0�}l���Hxh]�3tml�^P�l����̶��3�]����r��n5{�4p�j�[�l�
X��5D�Ss�x��FOq�П5.�gܷ�EÂg^��$,N��/PD���o��W�=��?㒛I�5�N`}�ߙk�.uzAM#�&���Z����^���a�;�\�$��w9K���H����4�G�,o:m�,q<D�[S��tTݧۃ��!r�J�0"�����"_������,�9�g�ց�H�e7�b��d�e1@L�un���|K�%5�TY�%�B�
+��F9����]����Pq������B���鶔"_��Ck��w�e�"ϙu� DG�J�j�w��OX*�Y4{"T>��Hɺܷ������G��N�\�dh�\U���_�<�9�)B��0�a^|T@�*>����po��eЌ�+�	�{���$�\�9X�,��	E��*���!�y�m���3{s�Lj.+V��^]����g�r�W)l�ҍY,Q������$��An�3��*G&�͢�5+��k�4��m�G�Ak��m�S�{B�(\�b��w:آ����b� �Ua�#�9hΏ�ۭ����W09�ӵ���5\Y�zI@���r�<������a^��#�-h���G}��@#90p?�ؠ�G��ٺI#)��"MK"V�1���ǔj�Ix�w`�"�C[ɘ�ۘ�69�t�\�Ǝ2�t�i9�$	�u�#������oe'Y�i�'b�<#�f2̭�e����	
����9@�[Z�;�;���	�!n Q�hܒ�C#��#���GJ�D�<nW�87�h�P�z���I�k���������M��Z�D�n!?N�q�g}Z��@�B��%�>��5U7(>3�-'�L�*9�I��Fk?��w8ipV�4��6)�A��e���D��ޏ� �j p�Ba�
�h�9�I���Z^9����7P(���������^"�j���0�d_FiB��Ձ��=D&�p��>8݇z{H�KP�!Q��_XH7RyJ��� �<�g�����'k��4n�].\9�eT���L�JÙ|��,D�2�ѳ��W�_�n��[�Y�����u��yA��Z���Q4tN����i�W���Iy���M�cb�
�?:�;i����ߐ����sH�>�ݚ�,E�6R{��9�v4ҫ�4�G�?D.̛u�p��5��"�� )bO���"���~`�%���#4R�o؟�lF!:h8,��Xawn�-�zR'�8>�1����>za<��������NCh���$Lݴ��"��侉�����c)����^��QR�S�H~*��~��噓�-���N�Q$�Օ4�'�`!�C�J?U����`w:=�0�}�p:ƍ=3�	�{X��%�������z�vD�c�|�(U�L������h��_�p�{^SzO� �Ƽ�
u+��ތoG\�?ݪKY�0Լ�Ǌ��+S����*v��'����Q��!GR�$�������]Y�z�,���B�����8�ĕl�3)�%;�Pr�;.��� 8p�_*��#u#��v$="���v�e����e�{�8ʝG��W�ϸ��ܸ�AT�XTk~Tl��J+�_��GGȄ�22�"�\%A4~�?��=�H��� �/�X	~��XYZ ]`鰿_5��ǀ�U..o�9������"`�W��2)i>�l���\n)��b���n3n3&߱`��l&"�P%�.1��Jh����Lf-
-�G�����@�����D?�X�o�Ǆ���3)@(�4s�],��������I�M-�)��VK�y��[,n�KNU�3�JU�5�� -j����k�U��8�\�yV���N�����vQ�L� 0�b��� VX1���ϔj��~���,����&�)j��4������l���~���yj��3�k�\]�$�=l=��-
��x.*�p���Ñ��a����J�֨���_���Z���P	�w�E#DԶ�%`Կ��XN���^1I]�L��Iv�14�:�����N��'�/�N��6VW���d����N8uek.yK�H᜷D�\$wf�@&�����I9%�̦���j��ᵊ�\��B��}̺a.&�*N��r"�s��䁃�]�+��l��2�v'�7Y���]��9:~�Fz�}�n2��~?H�juǖ�i��� =�����,�fr��HU�Zū��k�3����HB�m9WÅ�0Ĉ���6y�w[tR�2���ёj
�K
%�u(�V<\6:h�ǃs����|M[�P���K��:�;K��8�<{�����n��Hdu1�`��6�s���꟩T>ۡho%�#V�TD��x�
u�]@)�RO��(�|3ӑ���-2�"�_w \�zEюm��QEӐhp���z>�6���Ѕ��n�v0��x��ǌP����UZsX�`~�!�F�лy���i���^�n��p�S�&%xÄ��o��*2/v~��!*^<,���ЧU9|�Ѷ՚�(X����oܮ���D�Ed�׹�Ш��$v"އe;Y�W���
;�f��O,[��u��_���q�s���Q⦗��,!��/�Z��]��n�!��k�N��U,{I��6�%#�z���-�#+
�<����_X;�BJ˻����s�\b$�:��
,��5���\9�O<4�ܞ�)���/{\&hkr��	���*[��b"aǣ���l�����c4��ߊ���抹�L���d�����kQ�\m�\�/3_Y<�#6$f�B�D졌s_��(!�q�
�N~z��*��S����ǀ��ݒ}��u��������c�����Q�X�㚱"׬zϯ����h���p����^x5�͗��]t���o��+�*��4���C����
y�0�{w]0��{�5��c�Bx"N5yt!p�\ec�Wm[�!�����0��+�K��yn��Mz�s�z����(�
.;�������`�(�t�����$�݄=Q��;xJ|���n��Y_I�X����4p�UE
�ݿ�$�ca��T{���~��~�E�x�pI��~v3�Ա���?���J�S�ז�X�kWx�S�S��i�u��Y���p�^g�4����KDI7*EF�bW@۬X�>�ŏ뿕Xy6r�}ñ;�Kq�u��W��*���M�c��۾����
v�� ����t���ٯ(�2?��Y�Т����{�b�om�!'P8K�p��l��0р��\Fݔ� 5�r�j����f&����CO�2f�.��AodĪ�I��X/�MG�:	��|0v��6+�P�E�0�;���a�JQ7�!�^�s��|���^kHu<��O"ީD�R]A~\�_�Ji����g�!��Av��K	N�bm,�+hϯ�vm�ѽ��� ���46��2��֠BO{+s��:�-�i�y�s�ISݣw]����ʩDU���JD�4�.� ��>G��7'7����p"�K�[z�8l�8N�Dy����"��P.9��[���=�2���7
W�=���Ms�t�o�8d	)^�˪�^�5��n01`���O �q���RZ��)g�	��[���EG�z����&T�/���&��y=q~�ix���4N�s��_�.����oF�B�D�c���	���RK�nH�!d�Z�e��������h�n'�,��ЧP�����U~9�&V �$V����Ľ�99EiVwKm�+�:�_*+B�'������I[��J�>�Gf� A�k�:�L6+������3<2�m�
oµ��*CvC���,��捾���1��(�������K������mg�LB����K�����AK�Xh(5"���R]d�$�q�7�`E2G��i����R?�1�Ms�RĀjzU��C3w'�vWtɝfP7�/�v���S�x�*����s/�.�o��gQ���p�oa�T!��s�=�� ���^ddt�y�}�������X�]���17�Ĝ�|u��d�//��1�{_b����'�JDo/���аF�v��'��l��'{&�ʿ��(�.�݆���luE/cߪ�`��{v���WbF��1 ����d��iJ���rt) �`���t��̆�'���g����1?�N��I"��6�����Ap5��)�� �[��~����p�Z��h�X����V�a�
�(��CR�H���
��8*ܲ�`ŎsH��ʶJ�AT�F1������:����	)$]�����v��8Po��h��KU�F#��]���ݨ��]�Z���9hwF7���;Ws�e$���w������)�1��H)(�����`Jpk�*-�h��v]6hT���D�����H$�%�B����>�GDx��q�Ezq�@N,���
n�X�m�@��z &�\�Q��������l������9�R^`Q��~��0�"l���NY�i�%�5�X�[Sh�� �Ҿ)�%ob��BIc��6�ӂ=J
�������&�!��?��u���{��q��7|�X���M�
b`����}�Lw/i޵����}��䓀,�҅4�3��ܐ�ivyC	#�ɠp����B������Z�i@�V����n���K����u�����p�*;�M�iR�8��f%\������qs��U{Lv>�'|Ӵ��?���ID���&?3�Ⱥ���B��0)L��6�HV�SE�|v`�~���t`�������걾CC"I�7D�yN��Bӥ�ª��XB��Ε_�W�V5)�G*��26���bLy�����U'{����!���Ih{��!n���SF��DS�����/R��4yL��h�鱭������6�J���Vy�Y�mX�w�&��"�/?���q���V�x��[�xZ��ֽ <jK�EF��v%�;��u=Vo�K�RS�4>'�Hݻ�_�:���?��uɧ�+#I��ÿB�!��բ}3���U���������S�4�[��,��-J�-	�f�])��O�"�����:x����z\
�f.�G�*�X�*Y�(�*7����R<�)ۻ����f|U�c{�ߚ��ߋ�����*O:��L��h/�ӟ��Ba	��}\�>�)m6���9}%��_;Æe$�m.��v�r9����W�T�z���MT�ϗp�vm2�ί; ��=�:f�%��M4.��j��Ef9[�#�	W�x��yu\�^�k��t������;��q��; 4��sR5P�0��VZQ7/pJ�4��Ur�5e��J�DNj�	��;�xz_��R,�����
rR�>���9��� 4����*��'j,c�8� 與ȍ�w%g��!�կMDr�����
� ��:�ő������ѳ4w���|�\.�'͟���Gp�Ng���̎=у^d�C��fT�7���U���B�ƽ-�RR=1a�� ��7
Z�[ѓP[�4Ȣ[h��;��qXې�]����x�#A֬���d��[zM�������r��r^�x���
�e
�,�nlTE�%�x=j�I��T�z���}����I-Z�Jf�b~2J���`�U��蝗!D�U�`zD��2��.��O�2O���wAy
%c�1{
��#��U^�Ö�=�ލ�L��Ӎ��|3�=��m�s�{�/w�ڮ�ķ���XJ�4����.������N~��+Քx7�>��4
��q�w�%�RB���9sX�-re)��{>[�<�킜���Y��3�pNbx$g����xrܚ�߾�D\�Gh����E�k(J�&WG�p	Uj��z8�R�J�Vr|����1�����T�_Ȥ�~qȈ�و++7��9�x��;1@fBTaօ�#�s=,���H���m-.R�X��'�R��{���3�������,�!�NV�2¥$+4\����g�Үڗ��)��CJh:	3ģB�y}0��28��*y�
�Hك�\QCi��}��O��@��(8�pE/��r��Z��A%G����,}�@vQ�^45*�sb3��K���!ee��4�j1���c��7$�B��QJ1t$+n\����^�ﳅ ��}��S�o˥��J�<Tv�n��y��Pomٺ�.W65����^��{\УV���\���d��Z���&�:�tSQ���#O���}-y���~��_DU�I�/} S�G�V4Iޛ��3�ϵ�Q���(U�����k�{)h�{\':]�?����g_��I>��M*1��8������|T�͂���<$��R/�Z�t<k��~ܲV?>`~�j�S���d���+���+�kU�������cz,���K8�._@kX�>��!bgk�Q)��?1��	xП��D��KWע��7<�	��n�z�����'m\ؤ�dys�#i.�~��u o���'�׵>���$f�^b8������8��?������/
pa :E5^�/9�Q����={���h�;$�cr׫Rl@Teg�}�W�'z5��%��]�z9O$(�4M�#q���������W� ���ĸ�E�%a�����@U�;�8�DR��t:��hG�x�@bg*Q�7�~B'�o���8&�K:'}�h%�x�?(�Lt=��|���a�Z�d�	�k��� �9P���%�TL��]>U�g�_٢}�)p����A�s�?����3�I��]��b+d3�}H���G*�X菛_ղ��,2�?�P��X���b��zT�V�0pLێ!s�W�ڈ((I;�v�ٲ����v�SH'6C��3��(�������yz��*]�JP7/πJr.�\����S_��@�xѲ3�׸�=���F�uW�?n�@������y�S2~@OP�~���I������a�W�a����K?6����R�5�t�JE�����1�{�d�Gq���5\�
��y�/����D.A�Q[��;���X=o����(�롏�}�ZߙKnM�,����n1�}0�}�N��Ej�Q�"n*/W.'Y9���=��ճL�k�n%TK^%R��(��' |�w��<�a
���L���s�=�:�Ri��D(��f�:�R�w���Gt܎[F��������B�:uҶ���߆������z�I�$o�.�~�t?O���F�*��x��̐�gb�k�ARW�\y�VL����,rr��󎉛_�.�k���}��	ԍ���=.����ߖaL���L�(���?�[pn��={�x���B�M7��\<�_D]�֧*�HN�̩! �kNş�5�j�$���m}���gk��p�Z��	
&g����9\$!��k���]s������_�3����(��݂p\<ƙ�s�+�|7}K�nlDnD�ԯ<Dڿ�-���Y��o�����n۽����@z[�.E���i��z#��޳V3��zv�*��,��{mw|���#�MĎ!�#��3@z�I�_�ġ�p��%�m.�`D;#Mώ�2�@~�87mH;J2��6�",��QTp��{��.��,\c��E;M:B?�
(q�i���fܕA��*�����^��:�S���]��|#��>��~h~�	,o�h�=i%��
nV5�p@dO.�x?u��[��gn\��A�ߘ4�fy�f�vW�PW?����e�(a{��^I�},�r	�b���w�������_�C=4�Tok�ˌ����C�2;#@��!�@b9N��b>����_�U;aJ�>����#7��AӎB�'�]7Y\jF����@i���f�%gV�,������j�l�G^"��0��W��r��;K����i��J
@k�C0M���i<�V��Z�z��y㬊u�Df����c���aW����6_k%�h�oQ����k/�U��ƹ�{�4TٶzȿA�(�v��ԟ
^����!��؟5�~�"6�dFg���va�,
c�Ѝ�c��S�.�e�xe.f(��y�)��_�лbbꯁ9��R�f�73� !TQ��&�Z	�{BQ��B�v=�2�T���):B���YWu&MWreR30 ld�e}䲅श�Bg���8�D5�d�� �jPBdn�I��s����Z��=ߏ*z�����Ga<xϸ:] f��Y��!�����y���/��`�cyZPI�4Ɨ����`S\W�h(!��qz�_�ޘ���3�!�f�<eVh7F|9!/��/�m�hf�#lx�hb�qdt�	��@w&��̓Hྒྷϱ��!H϶��g?Ɓ��ےJR�6[^��>q���r&?�D����VRC����'g�c%Ɉ~�FDD蠭�m>�>V�yf�3pvdW\�D�z��h���,���W���L���N��C҅����2�+l�Jn����]Q���>p�XB�	���=�; pI�p[�9�s�{�(��E�^!�
" x��Me`��u�OoTpr��\-���(B8��e�j�[�Gps7�q\T$$���t��Y���Yp���"R	�>�^���زb��Ҷ�E��Ƙ�$ 4�\���_���޵#Fݿ�|9�멽Y�R���ux���v��aE����aU�����b;�E����ŧ��^��7��IL�r���8�A`�t�A�z��O�o�G"��!F�~���O2��lC�8�<1���`�����tA�CL\��M�4��S��<<�٭��D筫;�,��w^�7ܗ+=��F���']k`0W$/�fJNS�V��P�t�6���\�ؽ�U���lM���MF�Jz�Kp�3�,Q哓q�TD��ȍ�9��Y3�u��뾱��$]\���M
���oۀ��{a�Q�wc,� 7gh�q��T��u�<�Q<N �Ȕ>	��O�\_A�3g��q׾����O*&���q�����R�<��;��p���X'�u�M*@�;��p��ֻm�av�Q���K��ۛg��K�!/�@���@��}[(���W�����=o���SiIu��X�"vg-�"c�9u��	QM����L�� ��Cb�q�da'�`܁�O��`��,�]'���,��#%#GUJh�o������8n^��3�4���Қ��8~n���_OwԳ��J+�8A]��,��Xp�p5/�%a��4c!D3����U�ͨ���z;��dj=/JG"��5eYwU�_C�\�E�h!Js�ǈΉn����Ӿ�2��/�M�
����Mt3M�wpI�v�Z��(�f�0p�ԜL=YQ/P)�*p�L돥w���U���
!Z:'se`�}�q���������
���<t�W��h��$�_7Y�/)�$�[��~��
'�^�{����erNq�7�粼|��"�b���~��5Gu����7'!���s����E��������"n��6�a��{��;۷�t(e�7��BoF�b]b�ι�͹��H $#�L]�����vHf���!�-�0���nA��W��%�q�[0&貮����Ǚ��Q()K`F'l��hD��&�~�	�d'��5��udM� 8�LW�ο������[5S�=���'�@R�nt�O�r':���!rN@Dh0s����Us��@{�V�,����j��6��7������#;�PIU��Oɐ�epLY�pUYX��uz��)g�gF�\Ȅ )��ʐ���W$��vн9n�$�\r��(�
jI�c��ƫ�1O��Sy�i�{��Q�n��%|]��Yмp��^�gk�ŴksR��_���Ć����&���o7��ҡ��!���]G����;Q�z�?����1��}��d4a#���?@�r�n*��L�$+�$:������{s���E�Ψ�0�g��\kU*�pq���:x�( @�5�4�זƚ���='
�*��H�Tĥ�.���-�������+2*�>��8$鑇��|�&�d�{����H�8l.tYR΍qd>oH�xks�C�`��ȵN�)wN�]�e���Tx�Y���}p��=ze|��!��0&�tߺN��uT�ӌ��h�ne�l@lyDOX��	�VT(��V\��H�/�5�޼��as��8�
��\ w� zn6� ��8}Oi2��ӪPɢ��3�Z��f8��`��?�󦨉HX*�ʑ�8��;����똏L�R7�~C�y���$B�}9+Y}�g��K�<Z�Z��+#S$A�9�#��|���FKv��s��7���b8|�@��h)J���H(�z#�	d�i�\��4V:�^�a9����=�q��*�%��ZF70�y�����G�Wx����)ȹ}���Q�7��<c�De�x��/
'0$xG��o���)3-|�����_Hii�y���Gj	�30�3�8��ϡT4ꯨ\rœ�b��o��2 ��>�?��-�� ��ޘ���[����U�Tx�(����j�t���~�LiV���U"�)�Yc]T�x��H��`��rŘ��֐�@"�V�z�~R2, v������>ܽM��[�`��X��O�ت �̩7%݉�7`��D��pW0Z��*�X���s�����f�"e���G]΀�$�W�D��!�_	��",���H�zx��!�5P��.y�5g�5j�����˶
y �W�P[W��yc2#kbl��L|`��(��P�([.C��d7�JW~k
�帙V����+��q2�wӔcJ��T�t��`�5�yd2Pނ��`/0j&u���i0����F�T|ʽnV�gY��+Zܷ����@�2�+=KzB��d�;�Z��L� 7<�2�3�H��Ez|y�m$6G���-Ñ&����Oxw��Cw	ج��bГ𱜼��-is��p���_���		^�+�7
��y5���`��)mrP��c���ww�R���}�zI쵩��ٟ$nF�!�6Ճ��#��>`�H2Gh�LE�����"�z���tUx|7n0��@����M�N���oMf��̮�7�N5�*vα˔{�"	�&�)[�N[��F��Ҽ� ׇ�(��˛����|YT{��W�MUҸ��|�����9�#Q�[����߻N�.�#��_�|�~cL�>7�0��!�%|i(���292-��/��u�2v}�5cV8.��]ɏc��q����~7���� irC9]�1��	a���h|Y��o��3��	�d����7o)��b�;�>��?�&j��4��S&>UPx�An.��9�s�$"�w��h��'�.?�A��Auੑ&��G��ݹ��r��ĠKXA%x��.�0N�6Cw�NQ���I�Ջ�@K��8�܈���j��3��v)�����@��?
�K6��ma �;�B�wCOl���e�&�?o|�[�q��C�����l�AP��E��7�k"��Ac֩<kSE��v��ݲ�f��.�0�ҊT���#��|BM���x7UD�!�{!UO\��tM`S�V�i���"��V,B��$�4�bm�@6�W+�J�~�w[[�֙��8�,	J�K�ή��!�KIW�ȗ�87� J�^�U���5V#�;��=%����b��{>
�T��	���:���\��Ø�Sfl��M��Bd��Lr�1��> �	��z�W>����-e{��UB���N��_���o�� �����ѐ'��\QT�A��=�7��YE��B�u5ٰ�1���y�X�o����-��@��}����׶�_;ܒ�΁��� �*5�
ݒ}���4t w*54
�t��N��L�f�k�j����!�ǻ20@�\Ǵw@99e7�_w��d5Q��R�Ew�j��[	F�C	���O��ᜍ����9���KO7����2i)�>\S�@�.�r�\�O��^&�ߣ'�1f]�`����h���>�����-���'������lc������*'~���Bd���fp������^q�v8�C��3U���2y�X� ���M5j׶�GJ��szѯ���[ޔ-N�A<i;�@=�t��VƯ0A\��œ��Btf�]�.A��j���0m��?�,n'���8L�詒��ןt��Bllh,i[K�:�o��m���{����~|P�N�3	��X?���DQ%_�[��6�yӷ�`y�
�:�.���Y�ۑ�j�x6k�U������µ�c��V��rׇ[�H�p�}���o�[��NS�~C�f��-�b[�mO���[1g�)���،�V՝���#1N�!�O^��Z_5u���?�m'Y�Sv��e��"^�w��9p�n�Ka��e��0d�[��Y�7��
X�e����/��v���g�P���)�s�O�_���m�|�����4PB�(�Ί6g�s���M��}f'��U�����f^�#��`{�ЛU��?�ʓ��x�֣O/�_Ƞ�UxM����o�H�f|��k�-R����C�~�$�"���p��d��[���-8�O�HN��J���Ey�ab1'xbx ��amj^y#�.������Z�O��S��Sͭ���M��R�����y�CR�2����A� K�6�f�eO ��� ��!I%�Kn���<�qګ�����up�n����mb��D��Owc���[{OHߔG�[�g��`\Z`�ߧq����?�,~�۝Q�~�ɷ�e�ٰ|�d�.��ұ��W�΍97�B���(���!��O&�x��fø�Ҍ�l��B�Nf\A[�����rv�0м�}�Aqp�Z�c��a�St8�B�Ho+�H#҃����bI�u&� b8HOm�2��i��6@���b�1n6�&���N4�l���1L��&uǮ�ʁ1;y] *<���g�#��"ĪB)N�� #�m�,���t�y�-���jCƾ�n�4%���݂��x�t�d7NsA���y�I�^��;q��V�����tA$hǫy|�#�.�����ny;�-��du�%����)��WH;M�^={"o�#�x�=����m<6-�Ɛ�ߠ~�z5������!`��w	S��^������UG���C �e� �R�d��]N"DK����� ~2<���k�Am���Mܽ�1��O"��(f���>G)�2G�
�$�u
d���+��zL�ƫ	�+�W�A�r@ԗw	���Y�2�N ��&��CB}	�<5����`���P�����F��+�M����hD��K�en~d���^�}���~�4�r�9}��'�L�U�4����$��֬V
��ZBX%
1;I�mNl�]��}=�h�?�)r<�x9�t����
���aǪ��D�^�e���_����[x��}�0mL��!�?e-z���nFj���� ����ݟ�g[/�Ӫ_�_�ؤ[�ļ�J�1ʧ2K��j*]�����*,��%�cc!�{�ۃ��#'�#p�&v�@�7P���݃K�r�b�Q���Ȑ����[o|��ʫ���h�|�����!"&�b�c�Ɍ'gÒ����_��|���r8C9�\�{Kt+^����Wb�����G0�e�I���u��q�l���B-����9U�+��E!*YHHq���'�!Λ@�կ��0���&y���<��N�B
|�j»���G�S�o��a��u��}��$YI�YE��c�.�ڋxk�n[ ��cd3��Ɣ�;`w�MrbVm�"�^+�mwC�5�\�9Ewm��u�t��]���