library IEEE;
use IEEE.std_logic_1164.all;

entity initialisation is
	port (
		largeur_grille, hauteur_grille : out std_logic_vector(31 downto 0);
		--h_position_du_curseur, v_position_du_curseur : out std_logic_vector(31 downto 0);
		mode_jeu : out std_logic;
		type_grille : out std_logic;
		select_affichage : out std_logic;
		pause : out std_logic;
		map_init : out  std_logic_vector(1405 downto 0)
	);
end entity initialisation;

architecture a of initialisation is
begin

largeur_grille <= x"00000026";
hauteur_grille <= x"00000025";
--h_position_du_curseur <= x"00000001";
--v_position_du_curseur <= x"00000001";
mode_jeu <= '0';
type_grille <= '0';
select_affichage <= '1';
map_init(1405 downto 988) <= "0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000001010000000000000000000000000110000001100000000000011000000000000010001000011000000000000110011000000001000001000110000000000000000110000000010001011000010100000000000000000000000100000100000001000000000000000000000000100010000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000";
map_init(987 downto 0) <= (others => '0');
pause <= '0';
end architecture a;

--639 downto 0 =>"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000110000001100000000000011000000000000000000000000000000000000000100010000110000000000001100000000000000000000000000001100000000100000100011000000000000000000000000000000000000000000110000000010001011000010100000000000000000000000000000000000000000000000001000001000000010000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000"
--"000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010100000000000000000000000110000001100000000000011000000000001000100001100000000000011110000000010000010001100000000000000110000000010001011000010100000000000000000000010000010000000100000000000000000000001000100000000000000000000000000000000110000000000000000000000